library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is
	port(
		MAX10_CLK1_50 : in std_logic;
		KEY : in std_logic_vector(1 downto 0);

		VGA_B : out std_logic_vector(3 downto 0);
		VGA_G : out std_logic_vector(3 downto 0);
		VGA_R : out std_logic_vector(3 downto 0);
		VGA_HS : out std_logic;
		VGA_VS : out std_logic
	);
end entity top;

architecture arch of top is
	signal clock : std_logic;
	signal locked_sig : std_logic;
	component VGA
	port(
		clk : in std_logic;
		rst : in std_logic;

		blue : out std_logic_vector(3 downto 0);
		green : out std_logic_vector(3 downto 0);
		red : out std_logic_vector(3 downto 0);
		vgaHS : out std_logic;
		vgaVS : out std_logic
	);
	end component;
	
	component pll
	PORT(
		areset : in std_logic;
		inclk0 : in std_logic;
		c0 : out std_logic;
		locked : out std_logic
	);
	end component;

	begin
	pll_inst : pll
	PORT MAP(	
		areset => not KEY(0),
		inclk0 => MAX10_CLK1_50,
		c0 => clock,
		locked => locked_sig
	);

	VGATOP : VGA
	PORT MAP(
		clk => clock,
		rst => not KEY(0),

		blue => VGA_B,
		green => VGA_G,
		red => VGA_R,
		vgaHS => VGA_HS,
		vgaVS => VGA_VS
	);
end architecture arch;