LIBRARY ieee;
USE ieee.std_logic_1164.all;

entity audio_ctrl IS
	port (
        clk         : in  std_logic; -- 50 MHz, 50Mhz / 8kHz = 6250
        rst         : in  std_logic; 

        chompy_appy : in  std_logic; 
        twisty_turn : in  std_logic; 
        ha_loser    : in  std_logic; 

        audio_out   : out std_logic_vector(7 downto 0) -- GPIO(7 downto 0); 
	);
end audio_ctrl;

architecture arch OF audio_ctrl is 

    constant sine_len : integer := 128;
    constant vwoop_len : integer := 2000; 
    constant liz_len : integer := 7636; 
    constant womp_len : integer := 6431;


    type sine_table_t is array (0 to 127) of std_logic_vector(7 downto 0);
    
    type vwoop_table_t is array (0 to 1999)  of std_logic_vector(7 downto 0);
    type womp_table_t  is array (0 to 6430)  of std_logic_vector(7 downto 0);
    type liz_table_t is array (0 to 7636) of std_logic_vector(7 downto 0);

    signal lizLUT : liz_table_t := (
    0 => x"89",     1 => x"89",     2 => x"89",     3 => x"89",     4 => x"89",     5 => x"89",     6 => x"89",     7 => x"89", 
    8 => x"89",     9 => x"89",     10 => x"89",     11 => x"89",     12 => x"89",     13 => x"89",     14 => x"89",     15 => x"89", 
    16 => x"89",     17 => x"89",     18 => x"89",     19 => x"89",     20 => x"89",     21 => x"89",     22 => x"89",     23 => x"89", 
    24 => x"89",     25 => x"89",     26 => x"89",     27 => x"89",     28 => x"89",     29 => x"89",     30 => x"89",     31 => x"89", 
    32 => x"89",     33 => x"89",     34 => x"89",     35 => x"89",     36 => x"89",     37 => x"89",     38 => x"89",     39 => x"89", 
    40 => x"89",     41 => x"89",     42 => x"89",     43 => x"89",     44 => x"89",     45 => x"88",     46 => x"89",     47 => x"89", 
    48 => x"89",     49 => x"89",     50 => x"89",     51 => x"89",     52 => x"89",     53 => x"89",     54 => x"89",     55 => x"89", 
    56 => x"89",     57 => x"89",     58 => x"89",     59 => x"89",     60 => x"89",     61 => x"8A",     62 => x"89",     63 => x"8A", 
    64 => x"89",     65 => x"89",     66 => x"89",     67 => x"89",     68 => x"89",     69 => x"89",     70 => x"89",     71 => x"89", 
    72 => x"89",     73 => x"89",     74 => x"89",     75 => x"89",     76 => x"89",     77 => x"89",     78 => x"89",     79 => x"89", 
    80 => x"89",     81 => x"89",     82 => x"89",     83 => x"89",     84 => x"89",     85 => x"89",     86 => x"89",     87 => x"89", 
    88 => x"89",     89 => x"89",     90 => x"89",     91 => x"89",     92 => x"89",     93 => x"89",     94 => x"89",     95 => x"89", 
    96 => x"89",     97 => x"89",     98 => x"89",     99 => x"89",     100 => x"89",     101 => x"89",     102 => x"89",     103 => x"89", 
    104 => x"89",     105 => x"86",     106 => x"85",     107 => x"84",     108 => x"84",     109 => x"83",     110 => x"82",     111 => x"81", 
    112 => x"81",     113 => x"81",     114 => x"81",     115 => x"81",     116 => x"81",     117 => x"81",     118 => x"81",     119 => x"81", 
    120 => x"82",     121 => x"82",     122 => x"82",     123 => x"83",     124 => x"83",     125 => x"83",     126 => x"84",     127 => x"84", 
    128 => x"85",     129 => x"85",     130 => x"85",     131 => x"86",     132 => x"87",     133 => x"88",     134 => x"88",     135 => x"89", 
    136 => x"89",     137 => x"89",     138 => x"89",     139 => x"8A",     140 => x"8A",     141 => x"8A",     142 => x"8A",     143 => x"8A", 
    144 => x"8A",     145 => x"8A",     146 => x"8A",     147 => x"89",     148 => x"89",     149 => x"89",     150 => x"89",     151 => x"89", 
    152 => x"89",     153 => x"89",     154 => x"89",     155 => x"89",     156 => x"89",     157 => x"89",     158 => x"89",     159 => x"89", 
    160 => x"8A",     161 => x"8A",     162 => x"8A",     163 => x"8A",     164 => x"8A",     165 => x"8A",     166 => x"8A",     167 => x"8B", 
    168 => x"8B",     169 => x"8B",     170 => x"8B",     171 => x"8B",     172 => x"8C",     173 => x"8D",     174 => x"8D",     175 => x"8E", 
    176 => x"8E",     177 => x"8F",     178 => x"90",     179 => x"90",     180 => x"91",     181 => x"92",     182 => x"93",     183 => x"94", 
    184 => x"94",     185 => x"95",     186 => x"95",     187 => x"96",     188 => x"96",     189 => x"97",     190 => x"97",     191 => x"97", 
    192 => x"96",     193 => x"96",     194 => x"96",     195 => x"96",     196 => x"96",     197 => x"95",     198 => x"94",     199 => x"94", 
    200 => x"93",     201 => x"91",     202 => x"91",     203 => x"90",     204 => x"8F",     205 => x"8E",     206 => x"8D",     207 => x"8C", 
    208 => x"8C",     209 => x"8B",     210 => x"8A",     211 => x"8A",     212 => x"89",     213 => x"88",     214 => x"88",     215 => x"87", 
    216 => x"87",     217 => x"87",     218 => x"87",     219 => x"86",     220 => x"87",     221 => x"87",     222 => x"87",     223 => x"87", 
    224 => x"87",     225 => x"86",     226 => x"86",     227 => x"87",     228 => x"86",     229 => x"86",     230 => x"87",     231 => x"86", 
    232 => x"86",     233 => x"86",     234 => x"86",     235 => x"85",     236 => x"85",     237 => x"84",     238 => x"84",     239 => x"84", 
    240 => x"83",     241 => x"83",     242 => x"83",     243 => x"82",     244 => x"81",     245 => x"81",     246 => x"80",     247 => x"7F", 
    248 => x"7F",     249 => x"7E",     250 => x"7D",     251 => x"7D",     252 => x"7D",     253 => x"7C",     254 => x"7C",     255 => x"7C", 
    256 => x"7C",     257 => x"7C",     258 => x"7C",     259 => x"7C",     260 => x"7D",     261 => x"7D",     262 => x"7E",     263 => x"7E", 
    264 => x"7F",     265 => x"80",     266 => x"81",     267 => x"82",     268 => x"83",     269 => x"83",     270 => x"84",     271 => x"84", 
    272 => x"85",     273 => x"86",     274 => x"86",     275 => x"87",     276 => x"88",     277 => x"89",     278 => x"8A",     279 => x"8B", 
    280 => x"8B",     281 => x"8C",     282 => x"8D",     283 => x"8E",     284 => x"8F",     285 => x"8F",     286 => x"90",     287 => x"90", 
    288 => x"90",     289 => x"90",     290 => x"91",     291 => x"91",     292 => x"91",     293 => x"91",     294 => x"92",     295 => x"91", 
    296 => x"91",     297 => x"91",     298 => x"90",     299 => x"90",     300 => x"90",     301 => x"90",     302 => x"90",     303 => x"90", 
    304 => x"91",     305 => x"90",     306 => x"90",     307 => x"90",     308 => x"90",     309 => x"90",     310 => x"90",     311 => x"90", 
    312 => x"90",     313 => x"90",     314 => x"8F",     315 => x"8F",     316 => x"8F",     317 => x"8E",     318 => x"8E",     319 => x"8D", 
    320 => x"8E",     321 => x"8E",     322 => x"8D",     323 => x"8D",     324 => x"8C",     325 => x"8D",     326 => x"8D",     327 => x"8D", 
    328 => x"8D",     329 => x"8D",     330 => x"8D",     331 => x"8C",     332 => x"8B",     333 => x"8B",     334 => x"8A",     335 => x"8A", 
    336 => x"8A",     337 => x"8A",     338 => x"8A",     339 => x"89",     340 => x"89",     341 => x"87",     342 => x"86",     343 => x"85", 
    344 => x"84",     345 => x"83",     346 => x"83",     347 => x"83",     348 => x"83",     349 => x"82",     350 => x"81",     351 => x"81", 
    352 => x"80",     353 => x"80",     354 => x"80",     355 => x"80",     356 => x"80",     357 => x"81",     358 => x"81",     359 => x"81", 
    360 => x"81",     361 => x"81",     362 => x"82",     363 => x"82",     364 => x"83",     365 => x"83",     366 => x"84",     367 => x"85", 
    368 => x"85",     369 => x"85",     370 => x"85",     371 => x"86",     372 => x"86",     373 => x"88",     374 => x"88",     375 => x"89", 
    376 => x"89",     377 => x"88",     378 => x"89",     379 => x"88",     380 => x"89",     381 => x"89",     382 => x"89",     383 => x"89", 
    384 => x"8A",     385 => x"8A",     386 => x"89",     387 => x"89",     388 => x"89",     389 => x"88",     390 => x"88",     391 => x"88", 
    392 => x"88",     393 => x"89",     394 => x"89",     395 => x"89",     396 => x"89",     397 => x"89",     398 => x"88",     399 => x"88", 
    400 => x"88",     401 => x"88",     402 => x"88",     403 => x"88",     404 => x"89",     405 => x"89",     406 => x"89",     407 => x"89", 
    408 => x"89",     409 => x"89",     410 => x"8A",     411 => x"8A",     412 => x"8A",     413 => x"8A",     414 => x"8A",     415 => x"8B", 
    416 => x"8B",     417 => x"8C",     418 => x"8D",     419 => x"8E",     420 => x"8E",     421 => x"8E",     422 => x"8E",     423 => x"8F", 
    424 => x"8F",     425 => x"90",     426 => x"90",     427 => x"90",     428 => x"90",     429 => x"90",     430 => x"90",     431 => x"90", 
    432 => x"91",     433 => x"91",     434 => x"92",     435 => x"92",     436 => x"91",     437 => x"91",     438 => x"91",     439 => x"91", 
    440 => x"91",     441 => x"91",     442 => x"91",     443 => x"90",     444 => x"90",     445 => x"90",     446 => x"8F",     447 => x"8F", 
    448 => x"8E",     449 => x"8D",     450 => x"8D",     451 => x"8C",     452 => x"8C",     453 => x"8C",     454 => x"8C",     455 => x"8B", 
    456 => x"8B",     457 => x"8A",     458 => x"8A",     459 => x"89",     460 => x"89",     461 => x"89",     462 => x"88",     463 => x"88", 
    464 => x"88",     465 => x"88",     466 => x"88",     467 => x"87",     468 => x"86",     469 => x"86",     470 => x"86",     471 => x"85", 
    472 => x"85",     473 => x"85",     474 => x"84",     475 => x"84",     476 => x"82",     477 => x"81",     478 => x"81",     479 => x"80", 
    480 => x"80",     481 => x"80",     482 => x"80",     483 => x"7F",     484 => x"7F",     485 => x"7F",     486 => x"7E",     487 => x"7D", 
    488 => x"7D",     489 => x"7D",     490 => x"7E",     491 => x"7F",     492 => x"7F",     493 => x"80",     494 => x"80",     495 => x"80", 
    496 => x"80",     497 => x"81",     498 => x"82",     499 => x"83",     500 => x"84",     501 => x"85",     502 => x"86",     503 => x"86", 
    504 => x"87",     505 => x"87",     506 => x"87",     507 => x"88",     508 => x"89",     509 => x"8C",     510 => x"88",     511 => x"8A", 
    512 => x"8A",     513 => x"8D",     514 => x"8D",     515 => x"8B",     516 => x"88",     517 => x"8A",     518 => x"8F",     519 => x"92", 
    520 => x"92",     521 => x"88",     522 => x"86",     523 => x"8B",     524 => x"8F",     525 => x"91",     526 => x"8F",     527 => x"8F", 
    528 => x"8A",     529 => x"8A",     530 => x"8F",     531 => x"8E",     532 => x"91",     533 => x"8D",     534 => x"8E",     535 => x"8C", 
    536 => x"8D",     537 => x"91",     538 => x"8F",     539 => x"90",     540 => x"8E",     541 => x"8D",     542 => x"92",     543 => x"91", 
    544 => x"93",     545 => x"92",     546 => x"90",     547 => x"90",     548 => x"8D",     549 => x"8D",     550 => x"8E",     551 => x"91", 
    552 => x"96",     553 => x"93",     554 => x"90",     555 => x"8E",     556 => x"8D",     557 => x"8A",     558 => x"85",     559 => x"86", 
    560 => x"89",     561 => x"8B",     562 => x"89",     563 => x"89",     564 => x"89",     565 => x"87",     566 => x"85",     567 => x"85", 
    568 => x"81",     569 => x"81",     570 => x"85",     571 => x"87",     572 => x"89",     573 => x"89",     574 => x"84",     575 => x"83", 
    576 => x"82",     577 => x"84",     578 => x"82",     579 => x"82",     580 => x"85",     581 => x"87",     582 => x"88",     583 => x"85", 
    584 => x"83",     585 => x"82",     586 => x"82",     587 => x"82",     588 => x"83",     589 => x"84",     590 => x"85",     591 => x"88", 
    592 => x"8C",     593 => x"89",     594 => x"85",     595 => x"82",     596 => x"84",     597 => x"89",     598 => x"8A",     599 => x"8B", 
    600 => x"89",     601 => x"87",     602 => x"8A",     603 => x"8A",     604 => x"89",     605 => x"87",     606 => x"88",     607 => x"8A", 
    608 => x"8E",     609 => x"8F",     610 => x"8D",     611 => x"8D",     612 => x"8D",     613 => x"8E",     614 => x"8E",     615 => x"8D", 
    616 => x"8A",     617 => x"8B",     618 => x"8E",     619 => x"92",     620 => x"92",     621 => x"8E",     622 => x"8C",     623 => x"8E", 
    624 => x"90",     625 => x"90",     626 => x"8E",     627 => x"8C",     628 => x"8C",     629 => x"8C",     630 => x"8D",     631 => x"8E", 
    632 => x"8D",     633 => x"8E",     634 => x"8E",     635 => x"8F",     636 => x"8E",     637 => x"8C",     638 => x"8D",     639 => x"8E", 
    640 => x"8E",     641 => x"8E",     642 => x"8C",     643 => x"8C",     644 => x"8C",     645 => x"8D",     646 => x"8D",     647 => x"8B", 
    648 => x"8A",     649 => x"8A",     650 => x"8C",     651 => x"8C",     652 => x"8B",     653 => x"88",     654 => x"85",     655 => x"85", 
    656 => x"87",     657 => x"88",     658 => x"87",     659 => x"83",     660 => x"83",     661 => x"83",     662 => x"83",     663 => x"84", 
    664 => x"81",     665 => x"80",     666 => x"80",     667 => x"80",     668 => x"81",     669 => x"7F",     670 => x"7F",     671 => x"7E", 
    672 => x"7E",     673 => x"7F",     674 => x"7F",     675 => x"7F",     676 => x"80",     677 => x"80",     678 => x"80",     679 => x"7F", 
    680 => x"80",     681 => x"81",     682 => x"83",     683 => x"83",     684 => x"82",     685 => x"82",     686 => x"83",     687 => x"85", 
    688 => x"87",     689 => x"86",     690 => x"86",     691 => x"87",     692 => x"89",     693 => x"8A",     694 => x"8A",     695 => x"8B", 
    696 => x"8A",     697 => x"8A",     698 => x"8A",     699 => x"8C",     700 => x"8F",     701 => x"90",     702 => x"8E",     703 => x"8D", 
    704 => x"8E",     705 => x"90",     706 => x"93",     707 => x"94",     708 => x"93",     709 => x"91",     710 => x"91",     711 => x"93", 
    712 => x"93",     713 => x"92",     714 => x"92",     715 => x"91",     716 => x"90",     717 => x"8F",     718 => x"8E",     719 => x"8E", 
    720 => x"8F",     721 => x"90",     722 => x"8F",     723 => x"8D",     724 => x"8B",     725 => x"8C",     726 => x"8E",     727 => x"8F", 
    728 => x"8E",     729 => x"8C",     730 => x"8C",     731 => x"8C",     732 => x"8D",     733 => x"8E",     734 => x"8C",     735 => x"8C", 
    736 => x"8C",     737 => x"8C",     738 => x"8B",     739 => x"8A",     740 => x"8A",     741 => x"89",     742 => x"89",     743 => x"89", 
    744 => x"89",     745 => x"87",     746 => x"88",     747 => x"88",     748 => x"88",     749 => x"86",     750 => x"84",     751 => x"85", 
    752 => x"87",     753 => x"86",     754 => x"84",     755 => x"83",     756 => x"82",     757 => x"82",     758 => x"82",     759 => x"82", 
    760 => x"81",     761 => x"81",     762 => x"82",     763 => x"83",     764 => x"83",     765 => x"81",     766 => x"80",     767 => x"81", 
    768 => x"82",     769 => x"83",     770 => x"84",     771 => x"84",     772 => x"84",     773 => x"85",     774 => x"85",     775 => x"86", 
    776 => x"87",     777 => x"87",     778 => x"87",     779 => x"88",     780 => x"88",     781 => x"88",     782 => x"87",     783 => x"87", 
    784 => x"87",     785 => x"88",     786 => x"88",     787 => x"89",     788 => x"89",     789 => x"8A",     790 => x"8A",     791 => x"8A", 
    792 => x"8A",     793 => x"8A",     794 => x"8B",     795 => x"8C",     796 => x"8B",     797 => x"8B",     798 => x"8C",     799 => x"8C", 
    800 => x"8B",     801 => x"8B",     802 => x"8C",     803 => x"8D",     804 => x"8E",     805 => x"8D",     806 => x"8C",     807 => x"8C", 
    808 => x"8C",     809 => x"8C",     810 => x"8B",     811 => x"8A",     812 => x"8B",     813 => x"8B",     814 => x"8C",     815 => x"8D", 
    816 => x"8C",     817 => x"8B",     818 => x"8B",     819 => x"8B",     820 => x"8C",     821 => x"8B",     822 => x"8B",     823 => x"8B", 
    824 => x"8D",     825 => x"8D",     826 => x"8E",     827 => x"8D",     828 => x"8D",     829 => x"8D",     830 => x"8E",     831 => x"8F", 
    832 => x"8E",     833 => x"8F",     834 => x"8F",     835 => x"91",     836 => x"91",     837 => x"91",     838 => x"91",     839 => x"91", 
    840 => x"90",     841 => x"90",     842 => x"8F",     843 => x"8E",     844 => x"8E",     845 => x"8E",     846 => x"8E",     847 => x"8D", 
    848 => x"8D",     849 => x"8C",     850 => x"8C",     851 => x"8C",     852 => x"8C",     853 => x"8C",     854 => x"8C",     855 => x"8C", 
    856 => x"8C",     857 => x"8C",     858 => x"8C",     859 => x"8B",     860 => x"8B",     861 => x"8B",     862 => x"8B",     863 => x"8B", 
    864 => x"8B",     865 => x"8C",     866 => x"8B",     867 => x"8A",     868 => x"89",     869 => x"8A",     870 => x"8A",     871 => x"8A", 
    872 => x"89",     873 => x"88",     874 => x"88",     875 => x"87",     876 => x"87",     877 => x"87",     878 => x"85",     879 => x"85", 
    880 => x"84",     881 => x"84",     882 => x"83",     883 => x"83",     884 => x"83",     885 => x"83",     886 => x"83",     887 => x"83", 
    888 => x"82",     889 => x"82",     890 => x"81",     891 => x"81",     892 => x"81",     893 => x"82",     894 => x"82",     895 => x"82", 
    896 => x"82",     897 => x"81",     898 => x"81",     899 => x"80",     900 => x"80",     901 => x"81",     902 => x"81",     903 => x"82", 
    904 => x"82",     905 => x"81",     906 => x"80",     907 => x"7F",     908 => x"7F",     909 => x"80",     910 => x"81",     911 => x"81", 
    912 => x"81",     913 => x"81",     914 => x"81",     915 => x"81",     916 => x"82",     917 => x"82",     918 => x"83",     919 => x"83", 
    920 => x"84",     921 => x"85",     922 => x"86",     923 => x"87",     924 => x"87",     925 => x"87",     926 => x"87",     927 => x"88", 
    928 => x"89",     929 => x"89",     930 => x"8A",     931 => x"8B",     932 => x"8C",     933 => x"8C",     934 => x"8C",     935 => x"8C", 
    936 => x"8C",     937 => x"8C",     938 => x"8C",     939 => x"8C",     940 => x"8C",     941 => x"8C",     942 => x"8C",     943 => x"8C", 
    944 => x"8D",     945 => x"8C",     946 => x"8C",     947 => x"8C",     948 => x"8D",     949 => x"8E",     950 => x"8E",     951 => x"8E", 
    952 => x"8E",     953 => x"8E",     954 => x"8E",     955 => x"8D",     956 => x"8D",     957 => x"8D",     958 => x"8D",     959 => x"8E", 
    960 => x"90",     961 => x"90",     962 => x"90",     963 => x"90",     964 => x"8F",     965 => x"90",     966 => x"90",     967 => x"90", 
    968 => x"90",     969 => x"91",     970 => x"91",     971 => x"91",     972 => x"90",     973 => x"8F",     974 => x"8E",     975 => x"8E", 
    976 => x"8E",     977 => x"8F",     978 => x"8F",     979 => x"8E",     980 => x"8D",     981 => x"8D",     982 => x"8C",     983 => x"8C", 
    984 => x"8B",     985 => x"8B",     986 => x"8A",     987 => x"8A",     988 => x"8A",     989 => x"8A",     990 => x"8A",     991 => x"8A", 
    992 => x"8A",     993 => x"89",     994 => x"88",     995 => x"88",     996 => x"88",     997 => x"88",     998 => x"89",     999 => x"89", 
    1000 => x"88",     1001 => x"87",     1002 => x"87",     1003 => x"88",     1004 => x"88",     1005 => x"88",     1006 => x"88",     1007 => x"88", 
    1008 => x"89",     1009 => x"89",     1010 => x"89",     1011 => x"89",     1012 => x"89",     1013 => x"89",     1014 => x"8A",     1015 => x"8B", 
    1016 => x"8C",     1017 => x"8C",     1018 => x"8D",     1019 => x"8D",     1020 => x"8D",     1021 => x"8C",     1022 => x"8C",     1023 => x"8C", 
    1024 => x"8B",     1025 => x"8B",     1026 => x"8B",     1027 => x"8A",     1028 => x"8A",     1029 => x"8A",     1030 => x"89",     1031 => x"89", 
    1032 => x"89",     1033 => x"88",     1034 => x"88",     1035 => x"87",     1036 => x"87",     1037 => x"87",     1038 => x"87",     1039 => x"87", 
    1040 => x"86",     1041 => x"85",     1042 => x"85",     1043 => x"85",     1044 => x"85",     1045 => x"85",     1046 => x"85",     1047 => x"85", 
    1048 => x"86",     1049 => x"86",     1050 => x"85",     1051 => x"85",     1052 => x"84",     1053 => x"85",     1054 => x"86",     1055 => x"87", 
    1056 => x"87",     1057 => x"87",     1058 => x"87",     1059 => x"87",     1060 => x"86",     1061 => x"85",     1062 => x"85",     1063 => x"86", 
    1064 => x"86",     1065 => x"87",     1066 => x"87",     1067 => x"87",     1068 => x"86",     1069 => x"87",     1070 => x"87",     1071 => x"87", 
    1072 => x"87",     1073 => x"87",     1074 => x"88",     1075 => x"88",     1076 => x"89",     1077 => x"89",     1078 => x"88",     1079 => x"87", 
    1080 => x"86",     1081 => x"86",     1082 => x"86",     1083 => x"86",     1084 => x"86",     1085 => x"85",     1086 => x"84",     1087 => x"84", 
    1088 => x"84",     1089 => x"84",     1090 => x"83",     1091 => x"83",     1092 => x"82",     1093 => x"83",     1094 => x"84",     1095 => x"84", 
    1096 => x"85",     1097 => x"85",     1098 => x"85",     1099 => x"86",     1100 => x"87",     1101 => x"87",     1102 => x"88",     1103 => x"89", 
    1104 => x"8A",     1105 => x"8A",     1106 => x"8B",     1107 => x"8C",     1108 => x"8C",     1109 => x"8D",     1110 => x"8E",     1111 => x"90", 
    1112 => x"90",     1113 => x"90",     1114 => x"8F",     1115 => x"8E",     1116 => x"8E",     1117 => x"8F",     1118 => x"90",     1119 => x"90", 
    1120 => x"90",     1121 => x"90",     1122 => x"90",     1123 => x"90",     1124 => x"90",     1125 => x"91",     1126 => x"92",     1127 => x"93", 
    1128 => x"95",     1129 => x"96",     1130 => x"96",     1131 => x"97",     1132 => x"96",     1133 => x"96",     1134 => x"96",     1135 => x"97", 
    1136 => x"97",     1137 => x"98",     1138 => x"98",     1139 => x"98",     1140 => x"98",     1141 => x"98",     1142 => x"97",     1143 => x"96", 
    1144 => x"96",     1145 => x"95",     1146 => x"95",     1147 => x"94",     1148 => x"93",     1149 => x"92",     1150 => x"91",     1151 => x"91", 
    1152 => x"90",     1153 => x"8F",     1154 => x"8E",     1155 => x"8E",     1156 => x"8E",     1157 => x"8D",     1158 => x"8B",     1159 => x"8A", 
    1160 => x"88",     1161 => x"88",     1162 => x"87",     1163 => x"87",     1164 => x"86",     1165 => x"85",     1166 => x"83",     1167 => x"82", 
    1168 => x"80",     1169 => x"7F",     1170 => x"7D",     1171 => x"7D",     1172 => x"7D",     1173 => x"7D",     1174 => x"7C",     1175 => x"7C", 
    1176 => x"7B",     1177 => x"7B",     1178 => x"7B",     1179 => x"7B",     1180 => x"7B",     1181 => x"7C",     1182 => x"7C",     1183 => x"7C", 
    1184 => x"7C",     1185 => x"7C",     1186 => x"7C",     1187 => x"7B",     1188 => x"7B",     1189 => x"7A",     1190 => x"7B",     1191 => x"7B", 
    1192 => x"7B",     1193 => x"7A",     1194 => x"7A",     1195 => x"7A",     1196 => x"7A",     1197 => x"7A",     1198 => x"79",     1199 => x"7A", 
    1200 => x"7A",     1201 => x"7A",     1202 => x"7A",     1203 => x"7A",     1204 => x"7B",     1205 => x"7B",     1206 => x"7C",     1207 => x"7D", 
    1208 => x"7E",     1209 => x"7F",     1210 => x"80",     1211 => x"81",     1212 => x"81",     1213 => x"82",     1214 => x"83",     1215 => x"84", 
    1216 => x"85",     1217 => x"87",     1218 => x"88",     1219 => x"88",     1220 => x"89",     1221 => x"8B",     1222 => x"8B",     1223 => x"8C", 
    1224 => x"8D",     1225 => x"8D",     1226 => x"8E",     1227 => x"8F",     1228 => x"8F",     1229 => x"90",     1230 => x"90",     1231 => x"90", 
    1232 => x"90",     1233 => x"91",     1234 => x"91",     1235 => x"92",     1236 => x"92",     1237 => x"92",     1238 => x"93",     1239 => x"93", 
    1240 => x"94",     1241 => x"94",     1242 => x"95",     1243 => x"96",     1244 => x"97",     1245 => x"97",     1246 => x"98",     1247 => x"99", 
    1248 => x"99",     1249 => x"99",     1250 => x"99",     1251 => x"99",     1252 => x"99",     1253 => x"9A",     1254 => x"9A",     1255 => x"9A", 
    1256 => x"9A",     1257 => x"99",     1258 => x"98",     1259 => x"98",     1260 => x"98",     1261 => x"98",     1262 => x"97",     1263 => x"97", 
    1264 => x"97",     1265 => x"97",     1266 => x"96",     1267 => x"95",     1268 => x"94",     1269 => x"94",     1270 => x"93",     1271 => x"93", 
    1272 => x"92",     1273 => x"92",     1274 => x"91",     1275 => x"90",     1276 => x"8F",     1277 => x"8E",     1278 => x"8E",     1279 => x"8C", 
    1280 => x"8B",     1281 => x"8A",     1282 => x"89",     1283 => x"89",     1284 => x"89",     1285 => x"88",     1286 => x"88",     1287 => x"87", 
    1288 => x"87",     1289 => x"86",     1290 => x"85",     1291 => x"85",     1292 => x"84",     1293 => x"84",     1294 => x"84",     1295 => x"83", 
    1296 => x"83",     1297 => x"82",     1298 => x"82",     1299 => x"81",     1300 => x"81",     1301 => x"81",     1302 => x"81",     1303 => x"82", 
    1304 => x"81",     1305 => x"81",     1306 => x"80",     1307 => x"7F",     1308 => x"7F",     1309 => x"7F",     1310 => x"7E",     1311 => x"7E", 
    1312 => x"7D",     1313 => x"7D",     1314 => x"7D",     1315 => x"7C",     1316 => x"7B",     1317 => x"7B",     1318 => x"7B",     1319 => x"7B", 
    1320 => x"7A",     1321 => x"7A",     1322 => x"7A",     1323 => x"7A",     1324 => x"7B",     1325 => x"7B",     1326 => x"7B",     1327 => x"7B", 
    1328 => x"7C",     1329 => x"7D",     1330 => x"7E",     1331 => x"7F",     1332 => x"80",     1333 => x"81",     1334 => x"81",     1335 => x"82", 
    1336 => x"83",     1337 => x"84",     1338 => x"86",     1339 => x"86",     1340 => x"87",     1341 => x"89",     1342 => x"89",     1343 => x"8A", 
    1344 => x"8B",     1345 => x"8C",     1346 => x"8D",     1347 => x"8E",     1348 => x"8F",     1349 => x"90",     1350 => x"91",     1351 => x"92", 
    1352 => x"93",     1353 => x"93",     1354 => x"94",     1355 => x"95",     1356 => x"96",     1357 => x"96",     1358 => x"96",     1359 => x"96", 
    1360 => x"97",     1361 => x"96",     1362 => x"96",     1363 => x"96",     1364 => x"96",     1365 => x"96",     1366 => x"96",     1367 => x"95", 
    1368 => x"95",     1369 => x"94",     1370 => x"94",     1371 => x"93",     1372 => x"92",     1373 => x"92",     1374 => x"92",     1375 => x"91", 
    1376 => x"91",     1377 => x"90",     1378 => x"90",     1379 => x"90",     1380 => x"8F",     1381 => x"8E",     1382 => x"8D",     1383 => x"8D", 
    1384 => x"8C",     1385 => x"8C",     1386 => x"8B",     1387 => x"8A",     1388 => x"89",     1389 => x"89",     1390 => x"89",     1391 => x"89", 
    1392 => x"89",     1393 => x"89",     1394 => x"8A",     1395 => x"8A",     1396 => x"8B",     1397 => x"8B",     1398 => x"8B",     1399 => x"8B", 
    1400 => x"8C",     1401 => x"8C",     1402 => x"8C",     1403 => x"8C",     1404 => x"8C",     1405 => x"8C",     1406 => x"8C",     1407 => x"8B", 
    1408 => x"8B",     1409 => x"8A",     1410 => x"8A",     1411 => x"89",     1412 => x"89",     1413 => x"89",     1414 => x"88",     1415 => x"88", 
    1416 => x"87",     1417 => x"86",     1418 => x"85",     1419 => x"84",     1420 => x"84",     1421 => x"83",     1422 => x"82",     1423 => x"81", 
    1424 => x"81",     1425 => x"80",     1426 => x"80",     1427 => x"7F",     1428 => x"7F",     1429 => x"7F",     1430 => x"7F",     1431 => x"7F", 
    1432 => x"80",     1433 => x"80",     1434 => x"80",     1435 => x"81",     1436 => x"81",     1437 => x"82",     1438 => x"83",     1439 => x"83", 
    1440 => x"83",     1441 => x"84",     1442 => x"84",     1443 => x"84",     1444 => x"84",     1445 => x"84",     1446 => x"84",     1447 => x"85", 
    1448 => x"85",     1449 => x"84",     1450 => x"84",     1451 => x"83",     1452 => x"83",     1453 => x"83",     1454 => x"83",     1455 => x"82", 
    1456 => x"82",     1457 => x"82",     1458 => x"83",     1459 => x"83",     1460 => x"84",     1461 => x"84",     1462 => x"85",     1463 => x"85", 
    1464 => x"86",     1465 => x"86",     1466 => x"87",     1467 => x"88",     1468 => x"88",     1469 => x"88",     1470 => x"89",     1471 => x"89", 
    1472 => x"89",     1473 => x"89",     1474 => x"8A",     1475 => x"8A",     1476 => x"8A",     1477 => x"8A",     1478 => x"8A",     1479 => x"8A", 
    1480 => x"8A",     1481 => x"8A",     1482 => x"8A",     1483 => x"8A",     1484 => x"8A",     1485 => x"8A",     1486 => x"8A",     1487 => x"89", 
    1488 => x"89",     1489 => x"89",     1490 => x"89",     1491 => x"89",     1492 => x"89",     1493 => x"88",     1494 => x"89",     1495 => x"89", 
    1496 => x"89",     1497 => x"8A",     1498 => x"8A",     1499 => x"8B",     1500 => x"8C",     1501 => x"8C",     1502 => x"8D",     1503 => x"8E", 
    1504 => x"8F",     1505 => x"8F",     1506 => x"90",     1507 => x"91",     1508 => x"91",     1509 => x"91",     1510 => x"91",     1511 => x"91", 
    1512 => x"91",     1513 => x"91",     1514 => x"91",     1515 => x"90",     1516 => x"90",     1517 => x"90",     1518 => x"90",     1519 => x"90", 
    1520 => x"90",     1521 => x"8F",     1522 => x"8F",     1523 => x"8F",     1524 => x"8F",     1525 => x"90",     1526 => x"8F",     1527 => x"8F", 
    1528 => x"90",     1529 => x"91",     1530 => x"91",     1531 => x"92",     1532 => x"92",     1533 => x"92",     1534 => x"92",     1535 => x"92", 
    1536 => x"92",     1537 => x"92",     1538 => x"92",     1539 => x"91",     1540 => x"91",     1541 => x"91",     1542 => x"90",     1543 => x"90", 
    1544 => x"90",     1545 => x"90",     1546 => x"90",     1547 => x"90",     1548 => x"8F",     1549 => x"8F",     1550 => x"8F",     1551 => x"8E", 
    1552 => x"8E",     1553 => x"8E",     1554 => x"8E",     1555 => x"8E",     1556 => x"8E",     1557 => x"8D",     1558 => x"8D",     1559 => x"8C", 
    1560 => x"8B",     1561 => x"8B",     1562 => x"8A",     1563 => x"8A",     1564 => x"8A",     1565 => x"8A",     1566 => x"89",     1567 => x"88", 
    1568 => x"88",     1569 => x"87",     1570 => x"87",     1571 => x"85",     1572 => x"85",     1573 => x"84",     1574 => x"83",     1575 => x"82", 
    1576 => x"81",     1577 => x"80",     1578 => x"7F",     1579 => x"7E",     1580 => x"7D",     1581 => x"7C",     1582 => x"7B",     1583 => x"7A", 
    1584 => x"7A",     1585 => x"79",     1586 => x"79",     1587 => x"79",     1588 => x"79",     1589 => x"78",     1590 => x"78",     1591 => x"78", 
    1592 => x"79",     1593 => x"79",     1594 => x"79",     1595 => x"7A",     1596 => x"79",     1597 => x"7A",     1598 => x"7A",     1599 => x"7B", 
    1600 => x"7B",     1601 => x"7B",     1602 => x"7C",     1603 => x"7D",     1604 => x"7E",     1605 => x"7F",     1606 => x"80",     1607 => x"81", 
    1608 => x"82",     1609 => x"83",     1610 => x"84",     1611 => x"85",     1612 => x"87",     1613 => x"88",     1614 => x"89",     1615 => x"8A", 
    1616 => x"8A",     1617 => x"8A",     1618 => x"8B",     1619 => x"8B",     1620 => x"8B",     1621 => x"8B",     1622 => x"8A",     1623 => x"8A", 
    1624 => x"8A",     1625 => x"8A",     1626 => x"89",     1627 => x"88",     1628 => x"88",     1629 => x"88",     1630 => x"87",     1631 => x"87", 
    1632 => x"87",     1633 => x"88",     1634 => x"88",     1635 => x"89",     1636 => x"8A",     1637 => x"8B",     1638 => x"8B",     1639 => x"8B", 
    1640 => x"8D",     1641 => x"8E",     1642 => x"8E",     1643 => x"8E",     1644 => x"8E",     1645 => x"8F",     1646 => x"90",     1647 => x"90", 
    1648 => x"90",     1649 => x"91",     1650 => x"92",     1651 => x"92",     1652 => x"94",     1653 => x"93",     1654 => x"94",     1655 => x"95", 
    1656 => x"94",     1657 => x"95",     1658 => x"95",     1659 => x"95",     1660 => x"96",     1661 => x"97",     1662 => x"96",     1663 => x"97", 
    1664 => x"97",     1665 => x"97",     1666 => x"97",     1667 => x"96",     1668 => x"96",     1669 => x"96",     1670 => x"95",     1671 => x"95", 
    1672 => x"94",     1673 => x"95",     1674 => x"96",     1675 => x"95",     1676 => x"95",     1677 => x"95",     1678 => x"94",     1679 => x"94", 
    1680 => x"94",     1681 => x"93",     1682 => x"94",     1683 => x"94",     1684 => x"93",     1685 => x"93",     1686 => x"92",     1687 => x"91", 
    1688 => x"91",     1689 => x"90",     1690 => x"90",     1691 => x"8F",     1692 => x"8F",     1693 => x"8F",     1694 => x"8E",     1695 => x"8E", 
    1696 => x"8E",     1697 => x"8D",     1698 => x"8D",     1699 => x"8D",     1700 => x"8C",     1701 => x"8C",     1702 => x"8B",     1703 => x"8A", 
    1704 => x"8A",     1705 => x"89",     1706 => x"88",     1707 => x"87",     1708 => x"85",     1709 => x"84",     1710 => x"83",     1711 => x"82", 
    1712 => x"82",     1713 => x"81",     1714 => x"80",     1715 => x"80",     1716 => x"7E",     1717 => x"7D",     1718 => x"7C",     1719 => x"7B", 
    1720 => x"7B",     1721 => x"7C",     1722 => x"7A",     1723 => x"7B",     1724 => x"7B",     1725 => x"7B",     1726 => x"7B",     1727 => x"79", 
    1728 => x"7A",     1729 => x"7A",     1730 => x"7A",     1731 => x"7C",     1732 => x"7C",     1733 => x"7C",     1734 => x"7B",     1735 => x"7B", 
    1736 => x"7A",     1737 => x"7B",     1738 => x"7A",     1739 => x"7A",     1740 => x"7B",     1741 => x"7B",     1742 => x"7B",     1743 => x"7B", 
    1744 => x"7A",     1745 => x"7A",     1746 => x"7B",     1747 => x"7A",     1748 => x"7C",     1749 => x"7D",     1750 => x"7D",     1751 => x"7E", 
    1752 => x"80",     1753 => x"81",     1754 => x"82",     1755 => x"82",     1756 => x"83",     1757 => x"83",     1758 => x"84",     1759 => x"85", 
    1760 => x"86",     1761 => x"88",     1762 => x"89",     1763 => x"8A",     1764 => x"8B",     1765 => x"8C",     1766 => x"8D",     1767 => x"8E", 
    1768 => x"8F",     1769 => x"8F",     1770 => x"90",     1771 => x"91",     1772 => x"91",     1773 => x"92",     1774 => x"92",     1775 => x"92", 
    1776 => x"93",     1777 => x"92",     1778 => x"92",     1779 => x"92",     1780 => x"91",     1781 => x"90",     1782 => x"90",     1783 => x"8F", 
    1784 => x"8F",     1785 => x"8F",     1786 => x"90",     1787 => x"91",     1788 => x"91",     1789 => x"93",     1790 => x"91",     1791 => x"92", 
    1792 => x"93",     1793 => x"94",     1794 => x"93",     1795 => x"97",     1796 => x"8F",     1797 => x"9B",     1798 => x"95",     1799 => x"95", 
    1800 => x"9F",     1801 => x"8B",     1802 => x"9E",     1803 => x"91",     1804 => x"96",     1805 => x"9D",     1806 => x"92",     1807 => x"97", 
    1808 => x"91",     1809 => x"92",     1810 => x"95",     1811 => x"92",     1812 => x"96",     1813 => x"8C",     1814 => x"94",     1815 => x"8E", 
    1816 => x"90",     1817 => x"93",     1818 => x"88",     1819 => x"8F",     1820 => x"8A",     1821 => x"87",     1822 => x"90",     1823 => x"86", 
    1824 => x"8B",     1825 => x"8C",     1826 => x"85",     1827 => x"90",     1828 => x"88",     1829 => x"8C",     1830 => x"90",     1831 => x"8D", 
    1832 => x"91",     1833 => x"94",     1834 => x"90",     1835 => x"8D",     1836 => x"8C",     1837 => x"80",     1838 => x"85",     1839 => x"81", 
    1840 => x"7D",     1841 => x"84",     1842 => x"7D",     1843 => x"7F",     1844 => x"80",     1845 => x"7F",     1846 => x"82",     1847 => x"81", 
    1848 => x"81",     1849 => x"80",     1850 => x"81",     1851 => x"81",     1852 => x"80",     1853 => x"7D",     1854 => x"72",     1855 => x"70", 
    1856 => x"6B",     1857 => x"6A",     1858 => x"6F",     1859 => x"6E",     1860 => x"70",     1861 => x"79",     1862 => x"7A",     1863 => x"80", 
    1864 => x"85",     1865 => x"80",     1866 => x"8D",     1867 => x"8F",     1868 => x"96",     1869 => x"9F",     1870 => x"98",     1871 => x"9C", 
    1872 => x"97",     1873 => x"8F",     1874 => x"90",     1875 => x"85",     1876 => x"7E",     1877 => x"83",     1878 => x"72",     1879 => x"7B", 
    1880 => x"6F",     1881 => x"68",     1882 => x"73",     1883 => x"6B",     1884 => x"79",     1885 => x"82",     1886 => x"84",     1887 => x"94", 
    1888 => x"95",     1889 => x"A4",     1890 => x"A2",     1891 => x"A7",     1892 => x"A5",     1893 => x"A0",     1894 => x"A7",     1895 => x"9B", 
    1896 => x"99",     1897 => x"92",     1898 => x"82",     1899 => x"86",     1900 => x"7D",     1901 => x"7B",     1902 => x"81",     1903 => x"79", 
    1904 => x"84",     1905 => x"87",     1906 => x"8A",     1907 => x"93",     1908 => x"94",     1909 => x"9A",     1910 => x"A5",     1911 => x"A3", 
    1912 => x"AA",     1913 => x"A8",     1914 => x"A4",     1915 => x"9E",     1916 => x"94",     1917 => x"8B",     1918 => x"7E",     1919 => x"7D", 
    1920 => x"6D",     1921 => x"6D",     1922 => x"6E",     1923 => x"65",     1924 => x"74",     1925 => x"76",     1926 => x"7A",     1927 => x"8D", 
    1928 => x"8C",     1929 => x"A0",     1930 => x"A5",     1931 => x"A9",     1932 => x"AD",     1933 => x"A6",     1934 => x"A4",     1935 => x"9A", 
    1936 => x"91",     1937 => x"86",     1938 => x"74",     1939 => x"71",     1940 => x"67",     1941 => x"6F",     1942 => x"74",     1943 => x"74", 
    1944 => x"80",     1945 => x"7E",     1946 => x"8F",     1947 => x"9C",     1948 => x"A1",     1949 => x"B0",     1950 => x"B4",     1951 => x"B8", 
    1952 => x"C0",     1953 => x"B9",     1954 => x"B6",     1955 => x"AB",     1956 => x"99",     1957 => x"98",     1958 => x"86",     1959 => x"7B", 
    1960 => x"6A",     1961 => x"59",     1962 => x"5A",     1963 => x"50",     1964 => x"54",     1965 => x"5A",     1966 => x"5D",     1967 => x"71", 
    1968 => x"7C",     1969 => x"91",     1970 => x"9B",     1971 => x"A1",     1972 => x"B0",     1973 => x"AB",     1974 => x"B7",     1975 => x"AB", 
    1976 => x"A0",     1977 => x"97",     1978 => x"7F",     1979 => x"7D",     1980 => x"6C",     1981 => x"63",     1982 => x"61",     1983 => x"58", 
    1984 => x"61",     1985 => x"65",     1986 => x"6C",     1987 => x"7B",     1988 => x"7E",     1989 => x"93",     1990 => x"9F",     1991 => x"B0", 
    1992 => x"BC",     1993 => x"BB",     1994 => x"C3",     1995 => x"B1",     1996 => x"BB",     1997 => x"A1",     1998 => x"9E",     1999 => x"8E", 
    2000 => x"71",     2001 => x"77",     2002 => x"59",     2003 => x"56",     2004 => x"54",     2005 => x"44",     2006 => x"58",     2007 => x"58", 
    2008 => x"66",     2009 => x"76",     2010 => x"81",     2011 => x"91",     2012 => x"99",     2013 => x"A9",     2014 => x"A7",     2015 => x"AC", 
    2016 => x"A4",     2017 => x"94",     2018 => x"8F",     2019 => x"79",     2020 => x"71",     2021 => x"6D",     2022 => x"5C",     2023 => x"65", 
    2024 => x"60",     2025 => x"67",     2026 => x"76",     2027 => x"77",     2028 => x"85",     2029 => x"95",     2030 => x"9A",     2031 => x"B2", 
    2032 => x"B2",     2033 => x"BC",     2034 => x"BB",     2035 => x"BB",     2036 => x"B7",     2037 => x"B0",     2038 => x"AA",     2039 => x"91", 
    2040 => x"8C",     2041 => x"7A",     2042 => x"6D",     2043 => x"6B",     2044 => x"5A",     2045 => x"55",     2046 => x"5A",     2047 => x"5A", 
    2048 => x"6C",     2049 => x"76",     2050 => x"85",     2051 => x"91",     2052 => x"9D",     2053 => x"A8",     2054 => x"B1",     2055 => x"B1", 
    2056 => x"AD",     2057 => x"AA",     2058 => x"A0",     2059 => x"97",     2060 => x"93",     2061 => x"84",     2062 => x"7E",     2063 => x"7D", 
    2064 => x"74",     2065 => x"81",     2066 => x"7D",     2067 => x"7D",     2068 => x"8D",     2069 => x"89",     2070 => x"9E",     2071 => x"A5", 
    2072 => x"A7",     2073 => x"B2",     2074 => x"B2",     2075 => x"B4",     2076 => x"B8",     2077 => x"B2",     2078 => x"A7",     2079 => x"A4", 
    2080 => x"9A",     2081 => x"94",     2082 => x"8D",     2083 => x"80",     2084 => x"78",     2085 => x"76",     2086 => x"78",     2087 => x"7E", 
    2088 => x"7F",     2089 => x"88",     2090 => x"8B",     2091 => x"93",     2092 => x"9B",     2093 => x"9D",     2094 => x"9B",     2095 => x"93", 
    2096 => x"8D",     2097 => x"86",     2098 => x"7D",     2099 => x"77",     2100 => x"6D",     2101 => x"69",     2102 => x"6A",     2103 => x"64", 
    2104 => x"6D",     2105 => x"6F",     2106 => x"76",     2107 => x"87",     2108 => x"8D",     2109 => x"9B",     2110 => x"A4",     2111 => x"A7", 
    2112 => x"AA",     2113 => x"B2",     2114 => x"AA",     2115 => x"AD",     2116 => x"A7",     2117 => x"98",     2118 => x"99",     2119 => x"86", 
    2120 => x"7F",     2121 => x"77",     2122 => x"64",     2123 => x"60",     2124 => x"55",     2125 => x"57",     2126 => x"60",     2127 => x"5E", 
    2128 => x"67",     2129 => x"6B",     2130 => x"6F",     2131 => x"76",     2132 => x"79",     2133 => x"77",     2134 => x"75",     2135 => x"72", 
    2136 => x"69",     2137 => x"68",     2138 => x"66",     2139 => x"5E",     2140 => x"64",     2141 => x"62",     2142 => x"62",     2143 => x"6F", 
    2144 => x"6F",     2145 => x"7B",     2146 => x"87",     2147 => x"8C",     2148 => x"9A",     2149 => x"A0",     2150 => x"A0",     2151 => x"AB", 
    2152 => x"AE",     2153 => x"A9",     2154 => x"B2",     2155 => x"A3",     2156 => x"9F",     2157 => x"9D",     2158 => x"88",     2159 => x"8A", 
    2160 => x"7C",     2161 => x"6E",     2162 => x"73",     2163 => x"69",     2164 => x"70",     2165 => x"75",     2166 => x"7A",     2167 => x"81", 
    2168 => x"8D",     2169 => x"92",     2170 => x"95",     2171 => x"9D",     2172 => x"95",     2173 => x"93",     2174 => x"92",     2175 => x"83", 
    2176 => x"85",     2177 => x"7D",     2178 => x"72",     2179 => x"7B",     2180 => x"75",     2181 => x"78",     2182 => x"81",     2183 => x"81", 
    2184 => x"92",     2185 => x"9D",     2186 => x"A7",     2187 => x"B5",     2188 => x"BB",     2189 => x"BD",     2190 => x"CA",     2191 => x"CB", 
    2192 => x"CA",     2193 => x"CF",     2194 => x"BA",     2195 => x"BA",     2196 => x"B7",     2197 => x"A6",     2198 => x"A0",     2199 => x"87", 
    2200 => x"77",     2201 => x"76",     2202 => x"71",     2203 => x"72",     2204 => x"72",     2205 => x"7B",     2206 => x"81",     2207 => x"8D", 
    2208 => x"91",     2209 => x"91",     2210 => x"9D",     2211 => x"95",     2212 => x"95",     2213 => x"8E",     2214 => x"86",     2215 => x"81", 
    2216 => x"74",     2217 => x"71",     2218 => x"71",     2219 => x"71",     2220 => x"77",     2221 => x"82",     2222 => x"88",     2223 => x"90", 
    2224 => x"9A",     2225 => x"9C",     2226 => x"AE",     2227 => x"A1",     2228 => x"A6",     2229 => x"BB",     2230 => x"B6",     2231 => x"B1", 
    2232 => x"96",     2233 => x"9B",     2234 => x"AF",     2235 => x"A4",     2236 => x"9F",     2237 => x"99",     2238 => x"A1",     2239 => x"8B", 
    2240 => x"79",     2241 => x"7C",     2242 => x"71",     2243 => x"6F",     2244 => x"55",     2245 => x"58",     2246 => x"5A",     2247 => x"50", 
    2248 => x"5D",     2249 => x"58",     2250 => x"63",     2251 => x"6C",     2252 => x"66",     2253 => x"81",     2254 => x"8E",     2255 => x"8C", 
    2256 => x"86",     2257 => x"80",     2258 => x"8A",     2259 => x"7D",     2260 => x"68",     2261 => x"70",     2262 => x"82",     2263 => x"87", 
    2264 => x"73",     2265 => x"7B",     2266 => x"98",     2267 => x"8F",     2268 => x"73",     2269 => x"5F",     2270 => x"77",     2271 => x"8F", 
    2272 => x"7F",     2273 => x"89",     2274 => x"AE",     2275 => x"B8",     2276 => x"A3",     2277 => x"9E",     2278 => x"B7",     2279 => x"A6", 
    2280 => x"88",     2281 => x"82",     2282 => x"7C",     2283 => x"66",     2284 => x"4E",     2285 => x"4E",     2286 => x"57",     2287 => x"52", 
    2288 => x"4D",     2289 => x"5B",     2290 => x"7B",     2291 => x"8B",     2292 => x"8D",     2293 => x"8C",     2294 => x"87",     2295 => x"8F", 
    2296 => x"87",     2297 => x"77",     2298 => x"88",     2299 => x"8E",     2300 => x"8C",     2301 => x"9F",     2302 => x"AC",     2303 => x"B8", 
    2304 => x"91",     2305 => x"6B",     2306 => x"7A",     2307 => x"87",     2308 => x"95",     2309 => x"A2",     2310 => x"B8",     2311 => x"BB", 
    2312 => x"AA",     2313 => x"B8",     2314 => x"B5",     2315 => x"AB",     2316 => x"A7",     2317 => x"9A",     2318 => x"9C",     2319 => x"90", 
    2320 => x"8C",     2321 => x"84",     2322 => x"74",     2323 => x"7E",     2324 => x"7B",     2325 => x"76",     2326 => x"7E",     2327 => x"80", 
    2328 => x"7F",     2329 => x"75",     2330 => x"80",     2331 => x"91",     2332 => x"7E",     2333 => x"80",     2334 => x"99",     2335 => x"A8", 
    2336 => x"A9",     2337 => x"98",     2338 => x"99",     2339 => x"8F",     2340 => x"78",     2341 => x"71",     2342 => x"68",     2343 => x"75", 
    2344 => x"84",     2345 => x"95",     2346 => x"A8",     2347 => x"B7",     2348 => x"C0",     2349 => x"B1",     2350 => x"BB",     2351 => x"B8", 
    2352 => x"9D",     2353 => x"9E",     2354 => x"A6",     2355 => x"AE",     2356 => x"98",     2357 => x"8C",     2358 => x"96",     2359 => x"87", 
    2360 => x"84",     2361 => x"87",     2362 => x"89",     2363 => x"70",     2364 => x"59",     2365 => x"6C",     2366 => x"76",     2367 => x"66", 
    2368 => x"66",     2369 => x"89",     2370 => x"8D",     2371 => x"78",     2372 => x"7F",     2373 => x"83",     2374 => x"7C",     2375 => x"61", 
    2376 => x"5B",     2377 => x"6F",     2378 => x"6E",     2379 => x"74",     2380 => x"88",     2381 => x"A2",     2382 => x"A0",     2383 => x"97", 
    2384 => x"A8",     2385 => x"A2",     2386 => x"94",     2387 => x"8F",     2388 => x"99",     2389 => x"A3",     2390 => x"9D",     2391 => x"B3", 
    2392 => x"BA",     2393 => x"B1",     2394 => x"B5",     2395 => x"AB",     2396 => x"9C",     2397 => x"82",     2398 => x"81",     2399 => x"85", 
    2400 => x"57",     2401 => x"4D",     2402 => x"6B",     2403 => x"68",     2404 => x"58",     2405 => x"53",     2406 => x"64",     2407 => x"63", 
    2408 => x"40",     2409 => x"54",     2410 => x"6B",     2411 => x"5C",     2412 => x"58",     2413 => x"70",     2414 => x"8D",     2415 => x"75", 
    2416 => x"7C",     2417 => x"9B",     2418 => x"83",     2419 => x"76",     2420 => x"74",     2421 => x"88",     2422 => x"82",     2423 => x"7B", 
    2424 => x"AD",     2425 => x"AC",     2426 => x"B0",     2427 => x"D2",     2428 => x"D0",     2429 => x"BF",     2430 => x"B8",     2431 => x"C0", 
    2432 => x"A3",     2433 => x"84",     2434 => x"86",     2435 => x"89",     2436 => x"68",     2437 => x"48",     2438 => x"6C",     2439 => x"6C", 
    2440 => x"49",     2441 => x"59",     2442 => x"67",     2443 => x"5A",     2444 => x"4B",     2445 => x"62",     2446 => x"75",     2447 => x"6C", 
    2448 => x"7D",     2449 => x"8E",     2450 => x"88",     2451 => x"84",     2452 => x"93",     2453 => x"A1",     2454 => x"A1",     2455 => x"B1", 
    2456 => x"C8",     2457 => x"D0",     2458 => x"DF",     2459 => x"EE",     2460 => x"F5",     2461 => x"E5",     2462 => x"CB",     2463 => x"D9", 
    2464 => x"C7",     2465 => x"9A",     2466 => x"9D",     2467 => x"83",     2468 => x"6F",     2469 => x"71",     2470 => x"63",     2471 => x"70", 
    2472 => x"6B",     2473 => x"69",     2474 => x"78",     2475 => x"82",     2476 => x"85",     2477 => x"6A",     2478 => x"6F",     2479 => x"66", 
    2480 => x"4A",     2481 => x"4B",     2482 => x"49",     2483 => x"5F",     2484 => x"5A",     2485 => x"60",     2486 => x"8E",     2487 => x"95", 
    2488 => x"B3",     2489 => x"D2",     2490 => x"EC",     2491 => x"F8",     2492 => x"E0",     2493 => x"FF",     2494 => x"FC",     2495 => x"D2", 
    2496 => x"D4",     2497 => x"C5",     2498 => x"B6",     2499 => x"96",     2500 => x"7D",     2501 => x"7E",     2502 => x"64",     2503 => x"53", 
    2504 => x"58",     2505 => x"70",     2506 => x"7B",     2507 => x"77",     2508 => x"82",     2509 => x"6F",     2510 => x"5F",     2511 => x"5B", 
    2512 => x"4C",     2513 => x"4B",     2514 => x"3D",     2515 => x"4D",     2516 => x"63",     2517 => x"67",     2518 => x"8D",     2519 => x"A3", 
    2520 => x"A6",     2521 => x"A5",     2522 => x"BA",     2523 => x"DA",     2524 => x"C7",     2525 => x"C3",     2526 => x"CC",     2527 => x"CC", 
    2528 => x"C1",     2529 => x"9C",     2530 => x"95",     2531 => x"7F",     2532 => x"53",     2533 => x"49",     2534 => x"52",     2535 => x"5C", 
    2536 => x"51",     2537 => x"5D",     2538 => x"6F",     2539 => x"68",     2540 => x"67",     2541 => x"64",     2542 => x"6D",     2543 => x"60", 
    2544 => x"55",     2545 => x"73",     2546 => x"7C",     2547 => x"81",     2548 => x"94",     2549 => x"9C",     2550 => x"91",     2551 => x"94", 
    2552 => x"A3",     2553 => x"91",     2554 => x"8E",     2555 => x"A4",     2556 => x"B5",     2557 => x"B9",     2558 => x"B0",     2559 => x"B0", 
    2560 => x"9F",     2561 => x"6F",     2562 => x"4C",     2563 => x"4D",     2564 => x"3D",     2565 => x"2C",     2566 => x"43",     2567 => x"4D", 
    2568 => x"4A",     2569 => x"4B",     2570 => x"5E",     2571 => x"78",     2572 => x"78",     2573 => x"85",     2574 => x"9F",     2575 => x"B5", 
    2576 => x"C2",     2577 => x"D2",     2578 => x"D8",     2579 => x"BD",     2580 => x"B8",     2581 => x"AC",     2582 => x"90",     2583 => x"7D", 
    2584 => x"88",     2585 => x"AC",     2586 => x"9E",     2587 => x"A3",     2588 => x"BC",     2589 => x"A8",     2590 => x"8C",     2591 => x"7A", 
    2592 => x"83",     2593 => x"74",     2594 => x"63",     2595 => x"6E",     2596 => x"5F",     2597 => x"48",     2598 => x"34",     2599 => x"3C", 
    2600 => x"40",     2601 => x"37",     2602 => x"5E",     2603 => x"81",     2604 => x"9E",     2605 => x"C2",     2606 => x"D9",     2607 => x"E8", 
    2608 => x"E8",     2609 => x"E7",     2610 => x"E5",     2611 => x"CA",     2612 => x"BA",     2613 => x"D6",     2614 => x"DB",     2615 => x"C2", 
    2616 => x"C0",     2617 => x"BE",     2618 => x"A0",     2619 => x"7F",     2620 => x"79",     2621 => x"7A",     2622 => x"6A",     2623 => x"6A", 
    2624 => x"6A",     2625 => x"62",     2626 => x"55",     2627 => x"4C",     2628 => x"53",     2629 => x"46",     2630 => x"48",     2631 => x"61", 
    2632 => x"6F",     2633 => x"8B",     2634 => x"9E",     2635 => x"A0",     2636 => x"B5",     2637 => x"B6",     2638 => x"AC",     2639 => x"A0", 
    2640 => x"8A",     2641 => x"98",     2642 => x"A9",     2643 => x"A1",     2644 => x"A4",     2645 => x"AA",     2646 => x"A6",     2647 => x"93", 
    2648 => x"84",     2649 => x"87",     2650 => x"7B",     2651 => x"77",     2652 => x"7B",     2653 => x"71",     2654 => x"69",     2655 => x"57", 
    2656 => x"54",     2657 => x"55",     2658 => x"47",     2659 => x"5B",     2660 => x"72",     2661 => x"80",     2662 => x"97",     2663 => x"96", 
    2664 => x"9F",     2665 => x"A7",     2666 => x"97",     2667 => x"93",     2668 => x"7C",     2669 => x"78",     2670 => x"96",     2671 => x"93", 
    2672 => x"8E",     2673 => x"9D",     2674 => x"9B",     2675 => x"8B",     2676 => x"7D",     2677 => x"78",     2678 => x"6D",     2679 => x"61", 
    2680 => x"62",     2681 => x"63",     2682 => x"63",     2683 => x"51",     2684 => x"52",     2685 => x"62",     2686 => x"5F",     2687 => x"74", 
    2688 => x"8F",     2689 => x"A9",     2690 => x"CB",     2691 => x"CF",     2692 => x"DE",     2693 => x"F2",     2694 => x"DB",     2695 => x"C4", 
    2696 => x"AA",     2697 => x"96",     2698 => x"94",     2699 => x"7E",     2700 => x"75",     2701 => x"79",     2702 => x"6E",     2703 => x"6A", 
    2704 => x"66",     2705 => x"69",     2706 => x"66",     2707 => x"5E",     2708 => x"72",     2709 => x"71",     2710 => x"69",     2711 => x"69", 
    2712 => x"60",     2713 => x"66",     2714 => x"65",     2715 => x"73",     2716 => x"8E",     2717 => x"9F",     2718 => x"C4",     2719 => x"D6", 
    2720 => x"D9",     2721 => x"EA",     2722 => x"EC",     2723 => x"E2",     2724 => x"C9",     2725 => x"B9",     2726 => x"BE",     2727 => x"AA", 
    2728 => x"92",     2729 => x"88",     2730 => x"7E",     2731 => x"6C",     2732 => x"59",     2733 => x"5C",     2734 => x"5B",     2735 => x"52", 
    2736 => x"5A",     2737 => x"66",     2738 => x"72",     2739 => x"6E",     2740 => x"63",     2741 => x"6A",     2742 => x"64",     2743 => x"5D", 
    2744 => x"6C",     2745 => x"7F",     2746 => x"94",     2747 => x"9F",     2748 => x"A8",     2749 => x"BA",     2750 => x"C5",     2751 => x"C9", 
    2752 => x"C4",     2753 => x"BD",     2754 => x"C4",     2755 => x"C4",     2756 => x"AF",     2757 => x"9B",     2758 => x"92",     2759 => x"82", 
    2760 => x"63",     2761 => x"57",     2762 => x"5A",     2763 => x"4A",     2764 => x"3F",     2765 => x"43",     2766 => x"4C",     2767 => x"58", 
    2768 => x"55",     2769 => x"61",     2770 => x"79",     2771 => x"81",     2772 => x"96",     2773 => x"BA",     2774 => x"D5",     2775 => x"E5", 
    2776 => x"E6",     2777 => x"E8",     2778 => x"E9",     2779 => x"DB",     2780 => x"C9",     2781 => x"B6",     2782 => x"A3",     2783 => x"98", 
    2784 => x"8D",     2785 => x"76",     2786 => x"67",     2787 => x"60",     2788 => x"50",     2789 => x"41",     2790 => x"44",     2791 => x"4B", 
    2792 => x"4D",     2793 => x"4E",     2794 => x"53",     2795 => x"62",     2796 => x"64",     2797 => x"5E",     2798 => x"70",     2799 => x"77", 
    2800 => x"7A",     2801 => x"91",     2802 => x"A9",     2803 => x"C8",     2804 => x"D3",     2805 => x"D5",     2806 => x"EC",     2807 => x"F2", 
    2808 => x"F1",     2809 => x"EF",     2810 => x"E1",     2811 => x"D0",     2812 => x"BC",     2813 => x"A5",     2814 => x"84",     2815 => x"5E", 
    2816 => x"43",     2817 => x"2D",     2818 => x"12",     2819 => x"01",     2820 => x"03",     2821 => x"09",     2822 => x"0D",     2823 => x"19", 
    2824 => x"2D",     2825 => x"3B",     2826 => x"4B",     2827 => x"5B",     2828 => x"6E",     2829 => x"85",     2830 => x"96",     2831 => x"AB", 
    2832 => x"C1",     2833 => x"C9",     2834 => x"CD",     2835 => x"D3",     2836 => x"D7",     2837 => x"DD",     2838 => x"DE",     2839 => x"D6", 
    2840 => x"D1",     2841 => x"C8",     2842 => x"B7",     2843 => x"A6",     2844 => x"8F",     2845 => x"76",     2846 => x"60",     2847 => x"41", 
    2848 => x"27",     2849 => x"24",     2850 => x"21",     2851 => x"1D",     2852 => x"29",     2853 => x"34",     2854 => x"43",     2855 => x"4F", 
    2856 => x"5F",     2857 => x"7F",     2858 => x"91",     2859 => x"A0",     2860 => x"BA",     2861 => x"CB",     2862 => x"D4",     2863 => x"D7", 
    2864 => x"D8",     2865 => x"D8",     2866 => x"D4",     2867 => x"D0",     2868 => x"CC",     2869 => x"C8",     2870 => x"BF",     2871 => x"B6", 
    2872 => x"AE",     2873 => x"A5",     2874 => x"9C",     2875 => x"8C",     2876 => x"75",     2877 => x"61",     2878 => x"56",     2879 => x"55", 
    2880 => x"5B",     2881 => x"61",     2882 => x"6A",     2883 => x"74",     2884 => x"79",     2885 => x"86",     2886 => x"97",     2887 => x"A3", 
    2888 => x"AD",     2889 => x"B7",     2890 => x"C1",     2891 => x"C4",     2892 => x"C4",     2893 => x"C4",     2894 => x"C3",     2895 => x"BB", 
    2896 => x"AE",     2897 => x"A6",     2898 => x"A2",     2899 => x"94",     2900 => x"8B",     2901 => x"8B",     2902 => x"85",     2903 => x"7B", 
    2904 => x"6D",     2905 => x"62",     2906 => x"5B",     2907 => x"4F",     2908 => x"4E",     2909 => x"59",     2910 => x"61",     2911 => x"73", 
    2912 => x"81",     2913 => x"83",     2914 => x"8E",     2915 => x"9B",     2916 => x"A4",     2917 => x"A9",     2918 => x"AA",     2919 => x"B2", 
    2920 => x"B6",     2921 => x"AE",     2922 => x"A8",     2923 => x"A8",     2924 => x"9D",     2925 => x"92",     2926 => x"8D",     2927 => x"83", 
    2928 => x"77",     2929 => x"71",     2930 => x"72",     2931 => x"6C",     2932 => x"66",     2933 => x"66",     2934 => x"62",     2935 => x"55", 
    2936 => x"49",     2937 => x"4A",     2938 => x"55",     2939 => x"5B",     2940 => x"61",     2941 => x"70",     2942 => x"79",     2943 => x"81", 
    2944 => x"87",     2945 => x"8A",     2946 => x"92",     2947 => x"97",     2948 => x"9E",     2949 => x"A3",     2950 => x"A3",     2951 => x"A5", 
    2952 => x"A1",     2953 => x"9B",     2954 => x"94",     2955 => x"86",     2956 => x"79",     2957 => x"70",     2958 => x"6C",     2959 => x"67", 
    2960 => x"5D",     2961 => x"59",     2962 => x"5E",     2963 => x"62",     2964 => x"61",     2965 => x"65",     2966 => x"6A",     2967 => x"6E", 
    2968 => x"73",     2969 => x"7B",     2970 => x"83",     2971 => x"8B",     2972 => x"8F",     2973 => x"95",     2974 => x"98",     2975 => x"96", 
    2976 => x"94",     2977 => x"96",     2978 => x"98",     2979 => x"99",     2980 => x"99",     2981 => x"97",     2982 => x"94",     2983 => x"8E", 
    2984 => x"87",     2985 => x"84",     2986 => x"7E",     2987 => x"76",     2988 => x"74",     2989 => x"73",     2990 => x"6E",     2991 => x"6A", 
    2992 => x"69",     2993 => x"74",     2994 => x"80",     2995 => x"87",     2996 => x"8F",     2997 => x"97",     2998 => x"9E",     2999 => x"AB", 
    3000 => x"B6",     3001 => x"BB",     3002 => x"BA",     3003 => x"B7",     3004 => x"B3",     3005 => x"AD",     3006 => x"AA",     3007 => x"A8", 
    3008 => x"A4",     3009 => x"9E",     3010 => x"9D",     3011 => x"9F",     3012 => x"9D",     3013 => x"93",     3014 => x"8B",     3015 => x"85", 
    3016 => x"7E",     3017 => x"7A",     3018 => x"78",     3019 => x"72",     3020 => x"6E",     3021 => x"72",     3022 => x"7A",     3023 => x"80", 
    3024 => x"84",     3025 => x"8B",     3026 => x"93",     3027 => x"9B",     3028 => x"A3",     3029 => x"A9",     3030 => x"B1",     3031 => x"B6", 
    3032 => x"BB",     3033 => x"BB",     3034 => x"B9",     3035 => x"B9",     3036 => x"B6",     3037 => x"AD",     3038 => x"A8",     3039 => x"A0", 
    3040 => x"95",     3041 => x"87",     3042 => x"7D",     3043 => x"77",     3044 => x"71",     3045 => x"6C",     3046 => x"6E",     3047 => x"71", 
    3048 => x"6D",     3049 => x"6A",     3050 => x"6E",     3051 => x"71",     3052 => x"72",     3053 => x"73",     3054 => x"7A",     3055 => x"82", 
    3056 => x"86",     3057 => x"8B",     3058 => x"90",     3059 => x"92",     3060 => x"91",     3061 => x"91",     3062 => x"93",     3063 => x"97", 
    3064 => x"9B",     3065 => x"9E",     3066 => x"A0",     3067 => x"A3",     3068 => x"9F",     3069 => x"98",     3070 => x"8F",     3071 => x"83", 
    3072 => x"76",     3073 => x"6B",     3074 => x"62",     3075 => x"5E",     3076 => x"58",     3077 => x"55",     3078 => x"56",     3079 => x"5C", 
    3080 => x"5F",     3081 => x"63",     3082 => x"69",     3083 => x"70",     3084 => x"77",     3085 => x"7C",     3086 => x"84",     3087 => x"8A", 
    3088 => x"8F",     3089 => x"92",     3090 => x"93",     3091 => x"96",     3092 => x"99",     3093 => x"9C",     3094 => x"A0",     3095 => x"A0", 
    3096 => x"9F",     3097 => x"9C",     3098 => x"98",     3099 => x"92",     3100 => x"8A",     3101 => x"84",     3102 => x"7C",     3103 => x"74", 
    3104 => x"6E",     3105 => x"69",     3106 => x"64",     3107 => x"60",     3108 => x"5E",     3109 => x"5F",     3110 => x"5F",     3111 => x"60", 
    3112 => x"66",     3113 => x"70",     3114 => x"79",     3115 => x"80",     3116 => x"89",     3117 => x"93",     3118 => x"9C",     3119 => x"A6", 
    3120 => x"AC",     3121 => x"B7",     3122 => x"C3",     3123 => x"C6",     3124 => x"C9",     3125 => x"CA",     3126 => x"C7",     3127 => x"C0", 
    3128 => x"B8",     3129 => x"B0",     3130 => x"A6",     3131 => x"9C",     3132 => x"93",     3133 => x"8C",     3134 => x"84",     3135 => x"7D", 
    3136 => x"78",     3137 => x"72",     3138 => x"6A",     3139 => x"68",     3140 => x"67",     3141 => x"67",     3142 => x"6C",     3143 => x"72", 
    3144 => x"7B",     3145 => x"81",     3146 => x"87",     3147 => x"91",     3148 => x"99",     3149 => x"A3",     3150 => x"AF",     3151 => x"B9", 
    3152 => x"C0",     3153 => x"C2",     3154 => x"C3",     3155 => x"C2",     3156 => x"BC",     3157 => x"B4",     3158 => x"AB",     3159 => x"A0", 
    3160 => x"97",     3161 => x"8D",     3162 => x"83",     3163 => x"7D",     3164 => x"79",     3165 => x"73",     3166 => x"6C",     3167 => x"68", 
    3168 => x"6A",     3169 => x"68",     3170 => x"66",     3171 => x"68",     3172 => x"6C",     3173 => x"71",     3174 => x"73",     3175 => x"78", 
    3176 => x"80",     3177 => x"85",     3178 => x"8E",     3179 => x"99",     3180 => x"A2",     3181 => x"A8",     3182 => x"AB",     3183 => x"B0", 
    3184 => x"AF",     3185 => x"AA",     3186 => x"A4",     3187 => x"9C",     3188 => x"94",     3189 => x"8A",     3190 => x"83",     3191 => x"7C", 
    3192 => x"72",     3193 => x"6A",     3194 => x"61",     3195 => x"56",     3196 => x"50",     3197 => x"4A",     3198 => x"46",     3199 => x"47", 
    3200 => x"49",     3201 => x"4E",     3202 => x"55",     3203 => x"5D",     3204 => x"68",     3205 => x"72",     3206 => x"81",     3207 => x"91", 
    3208 => x"9F",     3209 => x"AD",     3210 => x"B9",     3211 => x"C2",     3212 => x"C9",     3213 => x"CB",     3214 => x"C9",     3215 => x"C1", 
    3216 => x"B8",     3217 => x"AE",     3218 => x"A1",     3219 => x"95",     3220 => x"8B",     3221 => x"7F",     3222 => x"73",     3223 => x"66", 
    3224 => x"5D",     3225 => x"55",     3226 => x"4E",     3227 => x"49",     3228 => x"48",     3229 => x"49",     3230 => x"4B",     3231 => x"4E", 
    3232 => x"53",     3233 => x"5A",     3234 => x"62",     3235 => x"6E",     3236 => x"7C",     3237 => x"89",     3238 => x"97",     3239 => x"A2", 
    3240 => x"AF",     3241 => x"B8",     3242 => x"BF",     3243 => x"C4",     3244 => x"C5",     3245 => x"C6",     3246 => x"C3",     3247 => x"BF", 
    3248 => x"BB",     3249 => x"B5",     3250 => x"AF",     3251 => x"A6",     3252 => x"9E",     3253 => x"96",     3254 => x"8D",     3255 => x"84", 
    3256 => x"7D",     3257 => x"76",     3258 => x"6E",     3259 => x"67",     3260 => x"63",     3261 => x"61",     3262 => x"60",     3263 => x"63", 
    3264 => x"68",     3265 => x"71",     3266 => x"7B",     3267 => x"86",     3268 => x"93",     3269 => x"9E",     3270 => x"A8",     3271 => x"B0", 
    3272 => x"B4",     3273 => x"B8",     3274 => x"B6",     3275 => x"B3",     3276 => x"AE",     3277 => x"A8",     3278 => x"A3",     3279 => x"9A", 
    3280 => x"93",     3281 => x"8D",     3282 => x"86",     3283 => x"81",     3284 => x"7C",     3285 => x"7A",     3286 => x"7C",     3287 => x"7F", 
    3288 => x"83",     3289 => x"88",     3290 => x"8D",     3291 => x"92",     3292 => x"97",     3293 => x"9B",     3294 => x"9E",     3295 => x"A2", 
    3296 => x"A7",     3297 => x"AB",     3298 => x"AA",     3299 => x"A9",     3300 => x"A8",     3301 => x"A7",     3302 => x"A3",     3303 => x"9C", 
    3304 => x"98",     3305 => x"92",     3306 => x"8C",     3307 => x"87",     3308 => x"82",     3309 => x"7D",     3310 => x"77",     3311 => x"70", 
    3312 => x"69",     3313 => x"62",     3314 => x"5E",     3315 => x"5D",     3316 => x"5D",     3317 => x"5E",     3318 => x"63",     3319 => x"69", 
    3320 => x"72",     3321 => x"7A",     3322 => x"81",     3323 => x"89",     3324 => x"90",     3325 => x"97",     3326 => x"9D",     3327 => x"A0", 
    3328 => x"A1",     3329 => x"A1",     3330 => x"9E",     3331 => x"9B",     3332 => x"97",     3333 => x"92",     3334 => x"8D",     3335 => x"89", 
    3336 => x"86",     3337 => x"82",     3338 => x"7F",     3339 => x"7C",     3340 => x"75",     3341 => x"6E",     3342 => x"67",     3343 => x"62", 
    3344 => x"5D",     3345 => x"5A",     3346 => x"58",     3347 => x"5C",     3348 => x"61",     3349 => x"65",     3350 => x"6B",     3351 => x"75", 
    3352 => x"7E",     3353 => x"87",     3354 => x"8F",     3355 => x"94",     3356 => x"99",     3357 => x"9A",     3358 => x"9A",     3359 => x"99", 
    3360 => x"94",     3361 => x"8F",     3362 => x"8A",     3363 => x"86",     3364 => x"83",     3365 => x"81",     3366 => x"82",     3367 => x"82", 
    3368 => x"82",     3369 => x"80",     3370 => x"7D",     3371 => x"7A",     3372 => x"78",     3373 => x"78",     3374 => x"77",     3375 => x"77", 
    3376 => x"7A",     3377 => x"7D",     3378 => x"81",     3379 => x"85",     3380 => x"8B",     3381 => x"93",     3382 => x"98",     3383 => x"9C", 
    3384 => x"A1",     3385 => x"A4",     3386 => x"A6",     3387 => x"A6",     3388 => x"A3",     3389 => x"A0",     3390 => x"9D",     3391 => x"99", 
    3392 => x"94",     3393 => x"92",     3394 => x"90",     3395 => x"8F",     3396 => x"8D",     3397 => x"88",     3398 => x"88",     3399 => x"87", 
    3400 => x"87",     3401 => x"88",     3402 => x"88",     3403 => x"8B",     3404 => x"8D",     3405 => x"90",     3406 => x"94",     3407 => x"98", 
    3408 => x"9D",     3409 => x"A2",     3410 => x"A7",     3411 => x"AC",     3412 => x"AE",     3413 => x"B1",     3414 => x"B1",     3415 => x"AF", 
    3416 => x"AB",     3417 => x"A7",     3418 => x"A3",     3419 => x"9B",     3420 => x"95",     3421 => x"90",     3422 => x"8B",     3423 => x"89", 
    3424 => x"85",     3425 => x"82",     3426 => x"80",     3427 => x"7C",     3428 => x"7B",     3429 => x"79",     3430 => x"78",     3431 => x"77", 
    3432 => x"77",     3433 => x"77",     3434 => x"79",     3435 => x"7A",     3436 => x"7F",     3437 => x"83",     3438 => x"87",     3439 => x"8C", 
    3440 => x"8F",     3441 => x"93",     3442 => x"96",     3443 => x"96",     3444 => x"95",     3445 => x"95",     3446 => x"92",     3447 => x"8F", 
    3448 => x"8E",     3449 => x"88",     3450 => x"85",     3451 => x"84",     3452 => x"82",     3453 => x"82",     3454 => x"7F",     3455 => x"7E", 
    3456 => x"80",     3457 => x"7C",     3458 => x"79",     3459 => x"78",     3460 => x"74",     3461 => x"70",     3462 => x"70",     3463 => x"71", 
    3464 => x"73",     3465 => x"75",     3466 => x"77",     3467 => x"7D",     3468 => x"81",     3469 => x"81",     3470 => x"84",     3471 => x"88", 
    3472 => x"87",     3473 => x"84",     3474 => x"7F",     3475 => x"7B",     3476 => x"78",     3477 => x"73",     3478 => x"70",     3479 => x"70", 
    3480 => x"70",     3481 => x"73",     3482 => x"75",     3483 => x"76",     3484 => x"7A",     3485 => x"7F",     3486 => x"82",     3487 => x"85", 
    3488 => x"88",     3489 => x"8E",     3490 => x"90",     3491 => x"8E",     3492 => x"8F",     3493 => x"93",     3494 => x"92",     3495 => x"92", 
    3496 => x"93",     3497 => x"96",     3498 => x"98",     3499 => x"96",     3500 => x"96",     3501 => x"94",     3502 => x"91",     3503 => x"8B", 
    3504 => x"86",     3505 => x"83",     3506 => x"7F",     3507 => x"7B",     3508 => x"79",     3509 => x"79",     3510 => x"7D",     3511 => x"7D", 
    3512 => x"7F",     3513 => x"85",     3514 => x"8B",     3515 => x"8E",     3516 => x"8D",     3517 => x"90",     3518 => x"96",     3519 => x"95", 
    3520 => x"93",     3521 => x"93",     3522 => x"94",     3523 => x"96",     3524 => x"93",     3525 => x"93",     3526 => x"97",     3527 => x"97", 
    3528 => x"95",     3529 => x"96",     3530 => x"99",     3531 => x"98",     3532 => x"97",     3533 => x"95",     3534 => x"9A",     3535 => x"99", 
    3536 => x"96",     3537 => x"97",     3538 => x"99",     3539 => x"95",     3540 => x"94",     3541 => x"95",     3542 => x"9C",     3543 => x"9E", 
    3544 => x"99",     3545 => x"97",     3546 => x"9B",     3547 => x"96",     3548 => x"93",     3549 => x"91",     3550 => x"8F",     3551 => x"90", 
    3552 => x"8C",     3553 => x"89",     3554 => x"8E",     3555 => x"8F",     3556 => x"8E",     3557 => x"90",     3558 => x"92",     3559 => x"96", 
    3560 => x"96",     3561 => x"93",     3562 => x"98",     3563 => x"99",     3564 => x"93",     3565 => x"91",     3566 => x"92",     3567 => x"92", 
    3568 => x"8D",     3569 => x"89",     3570 => x"89",     3571 => x"89",     3572 => x"82",     3573 => x"7C",     3574 => x"7A",     3575 => x"78", 
    3576 => x"71",     3577 => x"6D",     3578 => x"6C",     3579 => x"6C",     3580 => x"69",     3581 => x"6A",     3582 => x"6D",     3583 => x"72", 
    3584 => x"77",     3585 => x"7C",     3586 => x"82",     3587 => x"8A",     3588 => x"8E",     3589 => x"92",     3590 => x"97",     3591 => x"9C", 
    3592 => x"9F",     3593 => x"9A",     3594 => x"99",     3595 => x"9C",     3596 => x"99",     3597 => x"91",     3598 => x"8F",     3599 => x"8B", 
    3600 => x"84",     3601 => x"7B",     3602 => x"74",     3603 => x"73",     3604 => x"6C",     3605 => x"63",     3606 => x"61",     3607 => x"5F", 
    3608 => x"59",     3609 => x"57",     3610 => x"58",     3611 => x"5A",     3612 => x"5C",     3613 => x"5D",     3614 => x"68",     3615 => x"77", 
    3616 => x"7F",     3617 => x"8B",     3618 => x"98",     3619 => x"A3",     3620 => x"AB",     3621 => x"B0",     3622 => x"B4",     3623 => x"B8", 
    3624 => x"B6",     3625 => x"B2",     3626 => x"AC",     3627 => x"A0",     3628 => x"91",     3629 => x"84",     3630 => x"7A",     3631 => x"71", 
    3632 => x"67",     3633 => x"60",     3634 => x"5D",     3635 => x"5A",     3636 => x"59",     3637 => x"5D",     3638 => x"63",     3639 => x"6B", 
    3640 => x"70",     3641 => x"79",     3642 => x"86",     3643 => x"8D",     3644 => x"99",     3645 => x"A5",     3646 => x"A8",     3647 => x"AD", 
    3648 => x"B0",     3649 => x"B0",     3650 => x"B1",     3651 => x"AB",     3652 => x"A5",     3653 => x"A6",     3654 => x"A2",     3655 => x"99", 
    3656 => x"98",     3657 => x"94",     3658 => x"8D",     3659 => x"89",     3660 => x"85",     3661 => x"85",     3662 => x"82",     3663 => x"79", 
    3664 => x"79",     3665 => x"7A",     3666 => x"72",     3667 => x"70",     3668 => x"72",     3669 => x"76",     3670 => x"78",     3671 => x"7D", 
    3672 => x"87",     3673 => x"94",     3674 => x"9C",     3675 => x"A6",     3676 => x"B0",     3677 => x"B7",     3678 => x"BE",     3679 => x"BF", 
    3680 => x"BB",     3681 => x"B9",     3682 => x"B3",     3683 => x"A8",     3684 => x"9D",     3685 => x"91",     3686 => x"86",     3687 => x"78", 
    3688 => x"6B",     3689 => x"64",     3690 => x"60",     3691 => x"5D",     3692 => x"5D",     3693 => x"61",     3694 => x"66",     3695 => x"69", 
    3696 => x"72",     3697 => x"7F",     3698 => x"8A",     3699 => x"94",     3700 => x"9E",     3701 => x"A9",     3702 => x"B1",     3703 => x"B5", 
    3704 => x"B2",     3705 => x"B4",     3706 => x"B2",     3707 => x"A8",     3708 => x"A0",     3709 => x"A2",     3710 => x"9C",     3711 => x"8F", 
    3712 => x"85",     3713 => x"85",     3714 => x"8A",     3715 => x"85",     3716 => x"81",     3717 => x"8A",     3718 => x"91",     3719 => x"89", 
    3720 => x"88",     3721 => x"92",     3722 => x"92",     3723 => x"84",     3724 => x"82",     3725 => x"81",     3726 => x"79",     3727 => x"6D", 
    3728 => x"6D",     3729 => x"6F",     3730 => x"6D",     3731 => x"6B",     3732 => x"72",     3733 => x"7E",     3734 => x"87",     3735 => x"8B", 
    3736 => x"91",     3737 => x"99",     3738 => x"9D",     3739 => x"9A",     3740 => x"94",     3741 => x"91",     3742 => x"8C",     3743 => x"82", 
    3744 => x"74",     3745 => x"6B",     3746 => x"61",     3747 => x"57",     3748 => x"49",     3749 => x"45",     3750 => x"48",     3751 => x"4C", 
    3752 => x"51",     3753 => x"5A",     3754 => x"68",     3755 => x"78",     3756 => x"82",     3757 => x"8E",     3758 => x"9F",     3759 => x"AC", 
    3760 => x"B1",     3761 => x"BC",     3762 => x"C5",     3763 => x"C3",     3764 => x"BB",     3765 => x"B6",     3766 => x"AF",     3767 => x"9F", 
    3768 => x"8E",     3769 => x"85",     3770 => x"7B",     3771 => x"72",     3772 => x"75",     3773 => x"6D",     3774 => x"64",     3775 => x"63", 
    3776 => x"6C",     3777 => x"71",     3778 => x"78",     3779 => x"7F",     3780 => x"8F",     3781 => x"98",     3782 => x"97",     3783 => x"9E", 
    3784 => x"A6",     3785 => x"9A",     3786 => x"91",     3787 => x"93",     3788 => x"8A",     3789 => x"7F",     3790 => x"7A",     3791 => x"7A", 
    3792 => x"78",     3793 => x"76",     3794 => x"78",     3795 => x"80",     3796 => x"8C",     3797 => x"9C",     3798 => x"A3",     3799 => x"A8", 
    3800 => x"B0",     3801 => x"B5",     3802 => x"AD",     3803 => x"A8",     3804 => x"A7",     3805 => x"A2",     3806 => x"91",     3807 => x"7C", 
    3808 => x"76",     3809 => x"77",     3810 => x"69",     3811 => x"5F",     3812 => x"6B",     3813 => x"7B",     3814 => x"7F",     3815 => x"86", 
    3816 => x"9B",     3817 => x"B0",     3818 => x"B6",     3819 => x"C0",     3820 => x"D3",     3821 => x"DB",     3822 => x"D1",     3823 => x"CB", 
    3824 => x"D0",     3825 => x"C9",     3826 => x"B7",     3827 => x"A5",     3828 => x"9D",     3829 => x"93",     3830 => x"87",     3831 => x"7C", 
    3832 => x"78",     3833 => x"7D",     3834 => x"81",     3835 => x"7A",     3836 => x"7F",     3837 => x"96",     3838 => x"95",     3839 => x"81", 
    3840 => x"81",     3841 => x"96",     3842 => x"9C",     3843 => x"91",     3844 => x"91",     3845 => x"9D",     3846 => x"98",     3847 => x"7C", 
    3848 => x"73",     3849 => x"82",     3850 => x"77",     3851 => x"59",     3852 => x"54",     3853 => x"5A",     3854 => x"47",     3855 => x"33", 
    3856 => x"3C",     3857 => x"49",     3858 => x"46",     3859 => x"50",     3860 => x"6B",     3861 => x"7F",     3862 => x"92",     3863 => x"A4", 
    3864 => x"A8",     3865 => x"AD",     3866 => x"C1",     3867 => x"BD",     3868 => x"A0",     3869 => x"97",     3870 => x"9E",     3871 => x"86", 
    3872 => x"62",     3873 => x"5F",     3874 => x"68",     3875 => x"54",     3876 => x"43",     3877 => x"50",     3878 => x"64",     3879 => x"68", 
    3880 => x"6D",     3881 => x"7B",     3882 => x"8D",     3883 => x"95",     3884 => x"90",     3885 => x"8E",     3886 => x"99",     3887 => x"99", 
    3888 => x"88",     3889 => x"84",     3890 => x"89",     3891 => x"82",     3892 => x"74",     3893 => x"6E",     3894 => x"73",     3895 => x"76", 
    3896 => x"73",     3897 => x"74",     3898 => x"7C",     3899 => x"87",     3900 => x"88",     3901 => x"87",     3902 => x"92",     3903 => x"97", 
    3904 => x"92",     3905 => x"92",     3906 => x"94",     3907 => x"84",     3908 => x"76",     3909 => x"81",     3910 => x"8C",     3911 => x"7B", 
    3912 => x"64",     3913 => x"6B",     3914 => x"75",     3915 => x"68",     3916 => x"63",     3917 => x"77",     3918 => x"7D",     3919 => x"72", 
    3920 => x"74",     3921 => x"83",     3922 => x"89",     3923 => x"90",     3924 => x"9E",     3925 => x"AA",     3926 => x"B3",     3927 => x"C8", 
    3928 => x"D9",     3929 => x"DF",     3930 => x"E6",     3931 => x"EC",     3932 => x"DD",     3933 => x"CE",     3934 => x"D1",     3935 => x"CC", 
    3936 => x"A6",     3937 => x"8E",     3938 => x"9B",     3939 => x"97",     3940 => x"70",     3941 => x"6B",     3942 => x"87",     3943 => x"80", 
    3944 => x"61",     3945 => x"6F",     3946 => x"93",     3947 => x"97",     3948 => x"85",     3949 => x"8D",     3950 => x"9E",     3951 => x"9E", 
    3952 => x"94",     3953 => x"93",     3954 => x"96",     3955 => x"98",     3956 => x"94",     3957 => x"8F",     3958 => x"95",     3959 => x"9E", 
    3960 => x"98",     3961 => x"8D",     3962 => x"90",     3963 => x"96",     3964 => x"91",     3965 => x"86",     3966 => x"8A",     3967 => x"97", 
    3968 => x"98",     3969 => x"8B",     3970 => x"8C",     3971 => x"8F",     3972 => x"85",     3973 => x"7E",     3974 => x"85",     3975 => x"86", 
    3976 => x"83",     3977 => x"88",     3978 => x"90",     3979 => x"85",     3980 => x"6E",     3981 => x"73",     3982 => x"8D",     3983 => x"91", 
    3984 => x"83",     3985 => x"8B",     3986 => x"9D",     3987 => x"99",     3988 => x"90",     3989 => x"9D",     3990 => x"AD",     3991 => x"9F", 
    3992 => x"92",     3993 => x"9F",     3994 => x"A7",     3995 => x"9C",     3996 => x"98",     3997 => x"95",     3998 => x"84",     3999 => x"7B", 
    4000 => x"7F",     4001 => x"77",     4002 => x"64",     4003 => x"5D",     4004 => x"5E",     4005 => x"59",     4006 => x"58",     4007 => x"63", 
    4008 => x"62",     4009 => x"59",     4010 => x"6B",     4011 => x"86",     4012 => x"80",     4013 => x"72",     4014 => x"82",     4015 => x"91", 
    4016 => x"82",     4017 => x"6E",     4018 => x"72",     4019 => x"78",     4020 => x"6B",     4021 => x"59",     4022 => x"5A",     4023 => x"69", 
    4024 => x"6E",     4025 => x"65",     4026 => x"68",     4027 => x"79",     4028 => x"85",     4029 => x"8A",     4030 => x"8F",     4031 => x"93", 
    4032 => x"94",     4033 => x"94",     4034 => x"8E",     4035 => x"85",     4036 => x"82",     4037 => x"81",     4038 => x"7A",     4039 => x"74", 
    4040 => x"75",     4041 => x"7B",     4042 => x"79",     4043 => x"73",     4044 => x"76",     4045 => x"7C",     4046 => x"7C",     4047 => x"7C", 
    4048 => x"83",     4049 => x"88",     4050 => x"8B",     4051 => x"8D",     4052 => x"8C",     4053 => x"87",     4054 => x"94",     4055 => x"AB", 
    4056 => x"AC",     4057 => x"98",     4058 => x"9E",     4059 => x"B7",     4060 => x"BD",     4061 => x"AB",     4062 => x"AB",     4063 => x"B8", 
    4064 => x"AD",     4065 => x"8D",     4066 => x"88",     4067 => x"8D",     4068 => x"7B",     4069 => x"63",     4070 => x"5E",     4071 => x"60", 
    4072 => x"5B",     4073 => x"58",     4074 => x"5E",     4075 => x"64",     4076 => x"6A",     4077 => x"7C",     4078 => x"93",     4079 => x"A1", 
    4080 => x"AB",     4081 => x"BC",     4082 => x"C9",     4083 => x"CC",     4084 => x"D2",     4085 => x"D6",     4086 => x"C8",     4087 => x"B8", 
    4088 => x"BA",     4089 => x"B8",     4090 => x"9E",     4091 => x"8F",     4092 => x"97",     4093 => x"90",     4094 => x"71",     4095 => x"6A", 
    4096 => x"7D",     4097 => x"81",     4098 => x"76",     4099 => x"79",     4100 => x"83",     4101 => x"89",     4102 => x"8D",     4103 => x"90", 
    4104 => x"90",     4105 => x"99",     4106 => x"A4",     4107 => x"A6",     4108 => x"A2",     4109 => x"A9",     4110 => x"B1",     4111 => x"A7", 
    4112 => x"9B",     4113 => x"9D",     4114 => x"A1",     4115 => x"9B",     4116 => x"8F",     4117 => x"89",     4118 => x"90",     4119 => x"8F", 
    4120 => x"83",     4121 => x"80",     4122 => x"8A",     4123 => x"86",     4124 => x"79",     4125 => x"79",     4126 => x"85",     4127 => x"88", 
    4128 => x"84",     4129 => x"81",     4130 => x"86",     4131 => x"8C",     4132 => x"8A",     4133 => x"7A",     4134 => x"70",     4135 => x"7D", 
    4136 => x"8D",     4137 => x"80",     4138 => x"75",     4139 => x"8B",     4140 => x"98",     4141 => x"80",     4142 => x"7C",     4143 => x"96", 
    4144 => x"9B",     4145 => x"82",     4146 => x"7A",     4147 => x"82",     4148 => x"7B",     4149 => x"6C",     4150 => x"6C",     4151 => x"69", 
    4152 => x"55",     4153 => x"51",     4154 => x"65",     4155 => x"70",     4156 => x"69",     4157 => x"6D",     4158 => x"7F",     4159 => x"86", 
    4160 => x"83",     4161 => x"86",     4162 => x"8A",     4163 => x"8A",     4164 => x"8F",     4165 => x"91",     4166 => x"84",     4167 => x"77", 
    4168 => x"78",     4169 => x"78",     4170 => x"68",     4171 => x"5E",     4172 => x"6D",     4173 => x"77",     4174 => x"6C",     4175 => x"6A", 
    4176 => x"80",     4177 => x"8F",     4178 => x"89",     4179 => x"8A",     4180 => x"9A",     4181 => x"9F",     4182 => x"93",     4183 => x"8D", 
    4184 => x"91",     4185 => x"8F",     4186 => x"83",     4187 => x"7A",     4188 => x"75",     4189 => x"70",     4190 => x"71",     4191 => x"77", 
    4192 => x"7C",     4193 => x"81",     4194 => x"87",     4195 => x"8D",     4196 => x"91",     4197 => x"97",     4198 => x"9B",     4199 => x"9B", 
    4200 => x"99",     4201 => x"99",     4202 => x"98",     4203 => x"96",     4204 => x"97",     4205 => x"98",     4206 => x"93",     4207 => x"90", 
    4208 => x"93",     4209 => x"A0",     4210 => x"AC",     4211 => x"AD",     4212 => x"9F",     4213 => x"98",     4214 => x"9F",     4215 => x"A7", 
    4216 => x"9D",     4217 => x"95",     4218 => x"9C",     4219 => x"A0",     4220 => x"91",     4221 => x"8B",     4222 => x"95",     4223 => x"97", 
    4224 => x"88",     4225 => x"84",     4226 => x"8D",     4227 => x"8B",     4228 => x"79",     4229 => x"76",     4230 => x"7F",     4231 => x"82", 
    4232 => x"7C",     4233 => x"83",     4234 => x"94",     4235 => x"A0",     4236 => x"A5",     4237 => x"AC",     4238 => x"B2",     4239 => x"B2", 
    4240 => x"AF",     4241 => x"AD",     4242 => x"AE",     4243 => x"B1",     4244 => x"AC",     4245 => x"9C",     4246 => x"92",     4247 => x"93", 
    4248 => x"91",     4249 => x"7E",     4250 => x"73",     4251 => x"7F",     4252 => x"8C",     4253 => x"85",     4254 => x"7F",     4255 => x"8D", 
    4256 => x"9C",     4257 => x"97",     4258 => x"90",     4259 => x"96",     4260 => x"9A",     4261 => x"94",     4262 => x"92",     4263 => x"94", 
    4264 => x"8F",     4265 => x"7C",     4266 => x"6D",     4267 => x"67",     4268 => x"62",     4269 => x"59",     4270 => x"54",     4271 => x"57", 
    4272 => x"5F",     4273 => x"65",     4274 => x"6C",     4275 => x"74",     4276 => x"7B",     4277 => x"83",     4278 => x"8A",     4279 => x"90", 
    4280 => x"95",     4281 => x"98",     4282 => x"97",     4283 => x"97",     4284 => x"91",     4285 => x"84",     4286 => x"7A",     4287 => x"7B", 
    4288 => x"7F",     4289 => x"77",     4290 => x"68",     4291 => x"60",     4292 => x"64",     4293 => x"6E",     4294 => x"71",     4295 => x"6D", 
    4296 => x"6F",     4297 => x"76",     4298 => x"7C",     4299 => x"7E",     4300 => x"85",     4301 => x"8A",     4302 => x"86",     4303 => x"82", 
    4304 => x"83",     4305 => x"80",     4306 => x"75",     4307 => x"6E",     4308 => x"6D",     4309 => x"6A",     4310 => x"67",     4311 => x"6E", 
    4312 => x"7B",     4313 => x"80",     4314 => x"7F",     4315 => x"83",     4316 => x"8F",     4317 => x"96",     4318 => x"98",     4319 => x"9A", 
    4320 => x"A1",     4321 => x"A6",     4322 => x"A4",     4323 => x"A1",     4324 => x"A1",     4325 => x"9F",     4326 => x"99",     4327 => x"92", 
    4328 => x"8A",     4329 => x"88",     4330 => x"8B",     4331 => x"89",     4332 => x"7E",     4333 => x"79",     4334 => x"80",     4335 => x"84", 
    4336 => x"7B",     4337 => x"76",     4338 => x"80",     4339 => x"8F",     4340 => x"93",     4341 => x"92",     4342 => x"97",     4343 => x"9E", 
    4344 => x"9E",     4345 => x"9B",     4346 => x"9C",     4347 => x"9F",     4348 => x"A0",     4349 => x"9C",     4350 => x"97",     4351 => x"97", 
    4352 => x"9C",     4353 => x"9C",     4354 => x"95",     4355 => x"91",     4356 => x"96",     4357 => x"99",     4358 => x"94",     4359 => x"93", 
    4360 => x"9C",     4361 => x"A1",     4362 => x"9E",     4363 => x"9B",     4364 => x"A0",     4365 => x"A5",     4366 => x"A6",     4367 => x"A3", 
    4368 => x"A1",     4369 => x"A0",     4370 => x"9E",     4371 => x"96",     4372 => x"8E",     4373 => x"8E",     4374 => x"91",     4375 => x"90", 
    4376 => x"8B",     4377 => x"88",     4378 => x"87",     4379 => x"83",     4380 => x"7D",     4381 => x"7D",     4382 => x"7C",     4383 => x"78", 
    4384 => x"71",     4385 => x"6C",     4386 => x"62",     4387 => x"5A",     4388 => x"5C",     4389 => x"63",     4390 => x"62",     4391 => x"68", 
    4392 => x"79",     4393 => x"8A",     4394 => x"8F",     4395 => x"98",     4396 => x"A7",     4397 => x"B0",     4398 => x"B2",     4399 => x"B5", 
    4400 => x"B6",     4401 => x"B0",     4402 => x"AB",     4403 => x"A9",     4404 => x"9B",     4405 => x"86",     4406 => x"7E",     4407 => x"7C", 
    4408 => x"6D",     4409 => x"5B",     4410 => x"5D",     4411 => x"69",     4412 => x"69",     4413 => x"62",     4414 => x"67",     4415 => x"73", 
    4416 => x"77",     4417 => x"76",     4418 => x"7D",     4419 => x"87",     4420 => x"8B",     4421 => x"89",     4422 => x"86",     4423 => x"82", 
    4424 => x"81",     4425 => x"80",     4426 => x"78",     4427 => x"70",     4428 => x"74",     4429 => x"7B",     4430 => x"7C",     4431 => x"7D", 
    4432 => x"87",     4433 => x"90",     4434 => x"8E",     4435 => x"8D",     4436 => x"97",     4437 => x"9D",     4438 => x"98",     4439 => x"93", 
    4440 => x"95",     4441 => x"95",     4442 => x"8E",     4443 => x"89",     4444 => x"89",     4445 => x"85",     4446 => x"7E",     4447 => x"7F", 
    4448 => x"86",     4449 => x"89",     4450 => x"84",     4451 => x"84",     4452 => x"8E",     4453 => x"92",     4454 => x"87",     4455 => x"84", 
    4456 => x"92",     4457 => x"9E",     4458 => x"9A",     4459 => x"94",     4460 => x"9C",     4461 => x"9E",     4462 => x"93",     4463 => x"8D", 
    4464 => x"91",     4465 => x"8A",     4466 => x"79",     4467 => x"6E",     4468 => x"70",     4469 => x"6D",     4470 => x"65",     4471 => x"61", 
    4472 => x"65",     4473 => x"6D",     4474 => x"7A",     4475 => x"88",     4476 => x"98",     4477 => x"A9",     4478 => x"B6",     4479 => x"BA", 
    4480 => x"BD",     4481 => x"C6",     4482 => x"CA",     4483 => x"BF",     4484 => x"B6",     4485 => x"B8",     4486 => x"B0",     4487 => x"99", 
    4488 => x"88",     4489 => x"84",     4490 => x"7B",     4491 => x"68",     4492 => x"5F",     4493 => x"66",     4494 => x"6B",     4495 => x"68", 
    4496 => x"67",     4497 => x"70",     4498 => x"77",     4499 => x"78",     4500 => x"7A",     4501 => x"81",     4502 => x"8A",     4503 => x"91", 
    4504 => x"93",     4505 => x"93",     4506 => x"94",     4507 => x"95",     4508 => x"90",     4509 => x"86",     4510 => x"83",     4511 => x"8A", 
    4512 => x"8F",     4513 => x"8C",     4514 => x"8B",     4515 => x"92",     4516 => x"96",     4517 => x"93",     4518 => x"93",     4519 => x"98", 
    4520 => x"99",     4521 => x"97",     4522 => x"97",     4523 => x"98",     4524 => x"96",     4525 => x"93",     4526 => x"8E",     4527 => x"84", 
    4528 => x"7F",     4529 => x"7E",     4530 => x"7A",     4531 => x"73",     4532 => x"72",     4533 => x"76",     4534 => x"6F",     4535 => x"6A", 
    4536 => x"73",     4537 => x"79",     4538 => x"73",     4539 => x"72",     4540 => x"84",     4541 => x"8E",     4542 => x"88",     4543 => x"86", 
    4544 => x"8F",     4545 => x"90",     4546 => x"88",     4547 => x"88",     4548 => x"8A",     4549 => x"83",     4550 => x"7A",     4551 => x"7C", 
    4552 => x"7C",     4553 => x"76",     4554 => x"77",     4555 => x"7F",     4556 => x"84",     4557 => x"88",     4558 => x"93",     4559 => x"9E", 
    4560 => x"A2",     4561 => x"A8",     4562 => x"B0",     4563 => x"AF",     4564 => x"AA",     4565 => x"AA",     4566 => x"A7",     4567 => x"9A", 
    4568 => x"90",     4569 => x"8C",     4570 => x"7D",     4571 => x"68",     4572 => x"61",     4573 => x"61",     4574 => x"54",     4575 => x"44", 
    4576 => x"4B",     4577 => x"5A",     4578 => x"5C",     4579 => x"5A",     4580 => x"67",     4581 => x"78",     4582 => x"7F",     4583 => x"85", 
    4584 => x"93",     4585 => x"A2",     4586 => x"A7",     4587 => x"AA",     4588 => x"B2",     4589 => x"B7",     4590 => x"B6",     4591 => x"B0", 
    4592 => x"AA",     4593 => x"A5",     4594 => x"A3",     4595 => x"9E",     4596 => x"94",     4597 => x"8A",     4598 => x"86",     4599 => x"80", 
    4600 => x"75",     4601 => x"6F",     4602 => x"70",     4603 => x"6E",     4604 => x"68",     4605 => x"68",     4606 => x"71",     4607 => x"77", 
    4608 => x"78",     4609 => x"7D",     4610 => x"85",     4611 => x"89",     4612 => x"8C",     4613 => x"93",     4614 => x"9C",     4615 => x"A1", 
    4616 => x"A1",     4617 => x"A0",     4618 => x"9E",     4619 => x"9E",     4620 => x"9D",     4621 => x"9A",     4622 => x"97",     4623 => x"98", 
    4624 => x"9B",     4625 => x"96",     4626 => x"91",     4627 => x"95",     4628 => x"97",     4629 => x"91",     4630 => x"8B",     4631 => x"8F", 
    4632 => x"92",     4633 => x"8C",     4634 => x"85",     4635 => x"87",     4636 => x"8A",     4637 => x"8A",     4638 => x"8B",     4639 => x"8F", 
    4640 => x"94",     4641 => x"98",     4642 => x"9B",     4643 => x"9F",     4644 => x"A5",     4645 => x"AB",     4646 => x"AB",     4647 => x"A8", 
    4648 => x"A7",     4649 => x"A8",     4650 => x"A2",     4651 => x"9A",     4652 => x"95",     4653 => x"93",     4654 => x"8D",     4655 => x"86", 
    4656 => x"84",     4657 => x"84",     4658 => x"80",     4659 => x"7D",     4660 => x"7F",     4661 => x"82",     4662 => x"82",     4663 => x"81", 
    4664 => x"81",     4665 => x"83",     4666 => x"84",     4667 => x"85",     4668 => x"84",     4669 => x"83",     4670 => x"84",     4671 => x"85", 
    4672 => x"84",     4673 => x"85",     4674 => x"89",     4675 => x"8C",     4676 => x"89",     4677 => x"86",     4678 => x"86",     4679 => x"85", 
    4680 => x"7F",     4681 => x"7B",     4682 => x"79",     4683 => x"77",     4684 => x"74",     4685 => x"72",     4686 => x"72",     4687 => x"73", 
    4688 => x"74",     4689 => x"75",     4690 => x"7A",     4691 => x"7F",     4692 => x"85",     4693 => x"87",     4694 => x"88",     4695 => x"89", 
    4696 => x"8A",     4697 => x"87",     4698 => x"80",     4699 => x"7A",     4700 => x"79",     4701 => x"76",     4702 => x"6E",     4703 => x"69", 
    4704 => x"6A",     4705 => x"6D",     4706 => x"6A",     4707 => x"69",     4708 => x"6E",     4709 => x"76",     4710 => x"7B",     4711 => x"7D", 
    4712 => x"82",     4713 => x"87",     4714 => x"88",     4715 => x"88",     4716 => x"8A",     4717 => x"8A",     4718 => x"88",     4719 => x"87", 
    4720 => x"86",     4721 => x"84",     4722 => x"82",     4723 => x"83",     4724 => x"85",     4725 => x"87",     4726 => x"89",     4727 => x"8B", 
    4728 => x"8E",     4729 => x"90",     4730 => x"8F",     4731 => x"8E",     4732 => x"8F",     4733 => x"8F",     4734 => x"8D",     4735 => x"8B", 
    4736 => x"8A",     4737 => x"89",     4738 => x"88",     4739 => x"88",     4740 => x"8B",     4741 => x"8E",     4742 => x"90",     4743 => x"93", 
    4744 => x"96",     4745 => x"99",     4746 => x"9A",     4747 => x"99",     4748 => x"98",     4749 => x"96",     4750 => x"94",     4751 => x"93", 
    4752 => x"92",     4753 => x"92",     4754 => x"91",     4755 => x"91",     4756 => x"91",     4757 => x"92",     4758 => x"93",     4759 => x"93", 
    4760 => x"92",     4761 => x"91",     4762 => x"92",     4763 => x"93",     4764 => x"91",     4765 => x"91",     4766 => x"92",     4767 => x"90", 
    4768 => x"8E",     4769 => x"90",     4770 => x"91",     4771 => x"92",     4772 => x"96",     4773 => x"9D",     4774 => x"A2",     4775 => x"A5", 
    4776 => x"AA",     4777 => x"AF",     4778 => x"B1",     4779 => x"B1",     4780 => x"B0",     4781 => x"B0",     4782 => x"AD",     4783 => x"A8", 
    4784 => x"A2",     4785 => x"9D",     4786 => x"95",     4787 => x"8F",     4788 => x"8A",     4789 => x"87",     4790 => x"84",     4791 => x"82", 
    4792 => x"82",     4793 => x"84",     4794 => x"83",     4795 => x"81",     4796 => x"81",     4797 => x"83",     4798 => x"83",     4799 => x"82", 
    4800 => x"81",     4801 => x"83",     4802 => x"84",     4803 => x"83",     4804 => x"82",     4805 => x"84",     4806 => x"85",     4807 => x"86", 
    4808 => x"86",     4809 => x"89",     4810 => x"8B",     4811 => x"8B",     4812 => x"89",     4813 => x"87",     4814 => x"84",     4815 => x"80", 
    4816 => x"7C",     4817 => x"79",     4818 => x"78",     4819 => x"76",     4820 => x"76",     4821 => x"76",     4822 => x"76",     4823 => x"74", 
    4824 => x"72",     4825 => x"72",     4826 => x"71",     4827 => x"6F",     4828 => x"6F",     4829 => x"70",     4830 => x"70",     4831 => x"6E", 
    4832 => x"6E",     4833 => x"70",     4834 => x"71",     4835 => x"72",     4836 => x"74",     4837 => x"77",     4838 => x"79",     4839 => x"7A", 
    4840 => x"7B",     4841 => x"7B",     4842 => x"7A",     4843 => x"76",     4844 => x"73",     4845 => x"71",     4846 => x"6E",     4847 => x"6A", 
    4848 => x"66",     4849 => x"63",     4850 => x"61",     4851 => x"5F",     4852 => x"60",     4853 => x"64",     4854 => x"68",     4855 => x"6D", 
    4856 => x"73",     4857 => x"7C",     4858 => x"85",     4859 => x"8C",     4860 => x"92",     4861 => x"98",     4862 => x"9C",     4863 => x"9E", 
    4864 => x"9E",     4865 => x"9F",     4866 => x"9E",     4867 => x"9B",     4868 => x"98",     4869 => x"97",     4870 => x"95",     4871 => x"93", 
    4872 => x"91",     4873 => x"92",     4874 => x"94",     4875 => x"97",     4876 => x"99",     4877 => x"9A",     4878 => x"9C",     4879 => x"9E", 
    4880 => x"9D",     4881 => x"9D",     4882 => x"9F",     4883 => x"A0",     4884 => x"9D",     4885 => x"9A",     4886 => x"99",     4887 => x"99", 
    4888 => x"96",     4889 => x"95",     4890 => x"97",     4891 => x"9B",     4892 => x"9C",     4893 => x"9E",     4894 => x"A2",     4895 => x"A6", 
    4896 => x"A8",     4897 => x"AA",     4898 => x"AC",     4899 => x"AF",     4900 => x"B0",     4901 => x"AD",     4902 => x"A9",     4903 => x"A6", 
    4904 => x"A4",     4905 => x"A0",     4906 => x"9A",     4907 => x"96",     4908 => x"95",     4909 => x"93",     4910 => x"8F",     4911 => x"8B", 
    4912 => x"8B",     4913 => x"8C",     4914 => x"8C",     4915 => x"8B",     4916 => x"8C",     4917 => x"8D",     4918 => x"8B",     4919 => x"8A", 
    4920 => x"89",     4921 => x"88",     4922 => x"87",     4923 => x"87",     4924 => x"88",     4925 => x"8A",     4926 => x"8B",     4927 => x"8A", 
    4928 => x"87",     4929 => x"86",     4930 => x"88",     4931 => x"89",     4932 => x"87",     4933 => x"85",     4934 => x"85",     4935 => x"83", 
    4936 => x"81",     4937 => x"83",     4938 => x"88",     4939 => x"8A",     4940 => x"88",     4941 => x"86",     4942 => x"84",     4943 => x"82", 
    4944 => x"7F",     4945 => x"7B",     4946 => x"77",     4947 => x"75",     4948 => x"72",     4949 => x"6E",     4950 => x"6B",     4951 => x"6A", 
    4952 => x"69",     4953 => x"68",     4954 => x"69",     4955 => x"6C",     4956 => x"71",     4957 => x"74",     4958 => x"79",     4959 => x"7F", 
    4960 => x"84",     4961 => x"87",     4962 => x"88",     4963 => x"88",     4964 => x"89",     4965 => x"8A",     4966 => x"89",     4967 => x"87", 
    4968 => x"85",     4969 => x"84",     4970 => x"81",     4971 => x"7E",     4972 => x"7D",     4973 => x"7F",     4974 => x"80",     4975 => x"80", 
    4976 => x"81",     4977 => x"84",     4978 => x"87",     4979 => x"88",     4980 => x"88",     4981 => x"88",     4982 => x"88",     4983 => x"86", 
    4984 => x"85",     4985 => x"84",     4986 => x"83",     4987 => x"82",     4988 => x"82",     4989 => x"80",     4990 => x"7D",     4991 => x"7C", 
    4992 => x"7F",     4993 => x"81",     4994 => x"82",     4995 => x"84",     4996 => x"87",     4997 => x"89",     4998 => x"89",     4999 => x"8A", 
    5000 => x"8B",     5001 => x"8B",     5002 => x"8C",     5003 => x"8D",     5004 => x"8D",     5005 => x"8B",     5006 => x"89",     5007 => x"86", 
    5008 => x"83",     5009 => x"80",     5010 => x"80",     5011 => x"80",     5012 => x"81",     5013 => x"83",     5014 => x"86",     5015 => x"88", 
    5016 => x"8B",     5017 => x"8E",     5018 => x"92",     5019 => x"97",     5020 => x"9E",     5021 => x"A2",     5022 => x"A3",     5023 => x"A4", 
    5024 => x"A4",     5025 => x"A2",     5026 => x"9F",     5027 => x"9F",     5028 => x"9D",     5029 => x"98",     5030 => x"93",     5031 => x"91", 
    5032 => x"8D",     5033 => x"89",     5034 => x"86",     5035 => x"86",     5036 => x"85",     5037 => x"84",     5038 => x"85",     5039 => x"87", 
    5040 => x"8B",     5041 => x"8F",     5042 => x"93",     5043 => x"96",     5044 => x"99",     5045 => x"9B",     5046 => x"9C",     5047 => x"9F", 
    5048 => x"A0",     5049 => x"A1",     5050 => x"A1",     5051 => x"9F",     5052 => x"9C",     5053 => x"98",     5054 => x"94",     5055 => x"91", 
    5056 => x"8E",     5057 => x"8B",     5058 => x"89",     5059 => x"88",     5060 => x"88",     5061 => x"86",     5062 => x"85",     5063 => x"84", 
    5064 => x"84",     5065 => x"85",     5066 => x"85",     5067 => x"86",     5068 => x"87",     5069 => x"87",     5070 => x"86",     5071 => x"84", 
    5072 => x"82",     5073 => x"81",     5074 => x"81",     5075 => x"81",     5076 => x"81",     5077 => x"80",     5078 => x"80",     5079 => x"80", 
    5080 => x"7F",     5081 => x"7E",     5082 => x"7E",     5083 => x"7E",     5084 => x"7E",     5085 => x"7D",     5086 => x"7B",     5087 => x"7A", 
    5088 => x"7A",     5089 => x"7A",     5090 => x"79",     5091 => x"77",     5092 => x"76",     5093 => x"77",     5094 => x"78",     5095 => x"7A", 
    5096 => x"7E",     5097 => x"82",     5098 => x"84",     5099 => x"85",     5100 => x"86",     5101 => x"88",     5102 => x"8A",     5103 => x"8B", 
    5104 => x"8C",     5105 => x"8E",     5106 => x"8F",     5107 => x"8D",     5108 => x"8C",     5109 => x"8B",     5110 => x"8A",     5111 => x"88", 
    5112 => x"88",     5113 => x"88",     5114 => x"87",     5115 => x"85",     5116 => x"84",     5117 => x"83",     5118 => x"82",     5119 => x"82", 
    5120 => x"82",     5121 => x"83",     5122 => x"84",     5123 => x"85",     5124 => x"86",     5125 => x"87",     5126 => x"88",     5127 => x"89", 
    5128 => x"8A",     5129 => x"8B",     5130 => x"8B",     5131 => x"8C",     5132 => x"8C",     5133 => x"8D",     5134 => x"8D",     5135 => x"8E", 
    5136 => x"8F",     5137 => x"8F",     5138 => x"8E",     5139 => x"8E",     5140 => x"8F",     5141 => x"90",     5142 => x"90",     5143 => x"90", 
    5144 => x"90",     5145 => x"90",     5146 => x"8F",     5147 => x"8F",     5148 => x"8F",     5149 => x"8E",     5150 => x"8D",     5151 => x"8C", 
    5152 => x"8C",     5153 => x"8B",     5154 => x"8B",     5155 => x"8B",     5156 => x"8B",     5157 => x"8B",     5158 => x"8B",     5159 => x"8B", 
    5160 => x"8B",     5161 => x"8B",     5162 => x"8B",     5163 => x"8C",     5164 => x"8C",     5165 => x"8C",     5166 => x"8C",     5167 => x"8D", 
    5168 => x"8E",     5169 => x"8F",     5170 => x"8F",     5171 => x"90",     5172 => x"91",     5173 => x"92",     5174 => x"93",     5175 => x"93", 
    5176 => x"95",     5177 => x"97",     5178 => x"97",     5179 => x"97",     5180 => x"96",     5181 => x"97",     5182 => x"96",     5183 => x"95", 
    5184 => x"94",     5185 => x"94",     5186 => x"93",     5187 => x"91",     5188 => x"8F",     5189 => x"8E",     5190 => x"8C",     5191 => x"8A", 
    5192 => x"88",     5193 => x"89",     5194 => x"89",     5195 => x"89",     5196 => x"88",     5197 => x"89",     5198 => x"8B",     5199 => x"8C", 
    5200 => x"8D",     5201 => x"8E",     5202 => x"91",     5203 => x"92",     5204 => x"92",     5205 => x"94",     5206 => x"95",     5207 => x"97", 
    5208 => x"97",     5209 => x"96",     5210 => x"96",     5211 => x"96",     5212 => x"94",     5213 => x"92",     5214 => x"90",     5215 => x"8E", 
    5216 => x"8C",     5217 => x"88",     5218 => x"84",     5219 => x"81",     5220 => x"7E",     5221 => x"7B",     5222 => x"78",     5223 => x"75", 
    5224 => x"74",     5225 => x"73",     5226 => x"71",     5227 => x"70",     5228 => x"70",     5229 => x"71",     5230 => x"72",     5231 => x"72", 
    5232 => x"74",     5233 => x"76",     5234 => x"78",     5235 => x"79",     5236 => x"7B",     5237 => x"7E",     5238 => x"80",     5239 => x"82", 
    5240 => x"84",     5241 => x"86",     5242 => x"87",     5243 => x"87",     5244 => x"86",     5245 => x"85",     5246 => x"85",     5247 => x"83", 
    5248 => x"80",     5249 => x"7E",     5250 => x"7D",     5251 => x"7C",     5252 => x"7A",     5253 => x"78",     5254 => x"78",     5255 => x"79", 
    5256 => x"79",     5257 => x"7B",     5258 => x"7D",     5259 => x"7F",     5260 => x"81",     5261 => x"83",     5262 => x"85",     5263 => x"88", 
    5264 => x"89",     5265 => x"8A",     5266 => x"8A",     5267 => x"8B",     5268 => x"8B",     5269 => x"8A",     5270 => x"89",     5271 => x"89", 
    5272 => x"88",     5273 => x"88",     5274 => x"89",     5275 => x"89",     5276 => x"8A",     5277 => x"8A",     5278 => x"8B",     5279 => x"8B", 
    5280 => x"8C",     5281 => x"8C",     5282 => x"8C",     5283 => x"8C",     5284 => x"8C",     5285 => x"8C",     5286 => x"8C",     5287 => x"8C", 
    5288 => x"8C",     5289 => x"8C",     5290 => x"8D",     5291 => x"8E",     5292 => x"8F",     5293 => x"91",     5294 => x"93",     5295 => x"94", 
    5296 => x"95",     5297 => x"96",     5298 => x"97",     5299 => x"97",     5300 => x"97",     5301 => x"97",     5302 => x"97",     5303 => x"97", 
    5304 => x"98",     5305 => x"97",     5306 => x"97",     5307 => x"97",     5308 => x"97",     5309 => x"96",     5310 => x"96",     5311 => x"95", 
    5312 => x"95",     5313 => x"94",     5314 => x"92",     5315 => x"91",     5316 => x"90",     5317 => x"8F",     5318 => x"8E",     5319 => x"8E", 
    5320 => x"8F",     5321 => x"90",     5322 => x"91",     5323 => x"92",     5324 => x"92",     5325 => x"92",     5326 => x"93",     5327 => x"93", 
    5328 => x"92",     5329 => x"93",     5330 => x"93",     5331 => x"92",     5332 => x"90",     5333 => x"8E",     5334 => x"8E",     5335 => x"8D", 
    5336 => x"8D",     5337 => x"8D",     5338 => x"8F",     5339 => x"8F",     5340 => x"8F",     5341 => x"8E",     5342 => x"8D",     5343 => x"8C", 
    5344 => x"8B",     5345 => x"89",     5346 => x"88",     5347 => x"86",     5348 => x"84",     5349 => x"81",     5350 => x"7E",     5351 => x"7B", 
    5352 => x"78",     5353 => x"76",     5354 => x"75",     5355 => x"75",     5356 => x"76",     5357 => x"77",     5358 => x"78",     5359 => x"7A", 
    5360 => x"7C",     5361 => x"7E",     5362 => x"7F",     5363 => x"80",     5364 => x"82",     5365 => x"84",     5366 => x"85",     5367 => x"86", 
    5368 => x"87",     5369 => x"87",     5370 => x"86",     5371 => x"86",     5372 => x"87",     5373 => x"87",     5374 => x"88",     5375 => x"89", 
    5376 => x"89",     5377 => x"89",     5378 => x"88",     5379 => x"88",     5380 => x"87",     5381 => x"86",     5382 => x"85",     5383 => x"85", 
    5384 => x"85",     5385 => x"84",     5386 => x"83",     5387 => x"81",     5388 => x"81",     5389 => x"80",     5390 => x"80",     5391 => x"80", 
    5392 => x"81",     5393 => x"81",     5394 => x"81",     5395 => x"81",     5396 => x"80",     5397 => x"80",     5398 => x"7F",     5399 => x"80", 
    5400 => x"80",     5401 => x"81",     5402 => x"81",     5403 => x"82",     5404 => x"83",     5405 => x"83",     5406 => x"84",     5407 => x"84", 
    5408 => x"85",     5409 => x"86",     5410 => x"87",     5411 => x"89",     5412 => x"8A",     5413 => x"8C",     5414 => x"8D",     5415 => x"8F", 
    5416 => x"90",     5417 => x"92",     5418 => x"93",     5419 => x"95",     5420 => x"96",     5421 => x"98",     5422 => x"99",     5423 => x"9A", 
    5424 => x"9B",     5425 => x"9B",     5426 => x"9C",     5427 => x"9C",     5428 => x"9D",     5429 => x"9C",     5430 => x"9C",     5431 => x"9C", 
    5432 => x"9B",     5433 => x"99",     5434 => x"97",     5435 => x"95",     5436 => x"94",     5437 => x"93",     5438 => x"91",     5439 => x"90", 
    5440 => x"8F",     5441 => x"8E",     5442 => x"8C",     5443 => x"8A",     5444 => x"89",     5445 => x"88",     5446 => x"87",     5447 => x"87", 
    5448 => x"86",     5449 => x"86",     5450 => x"86",     5451 => x"85",     5452 => x"85",     5453 => x"86",     5454 => x"87",     5455 => x"88", 
    5456 => x"89",     5457 => x"8B",     5458 => x"8C",     5459 => x"8E",     5460 => x"8F",     5461 => x"8F",     5462 => x"90",     5463 => x"91", 
    5464 => x"92",     5465 => x"93",     5466 => x"94",     5467 => x"94",     5468 => x"94",     5469 => x"94",     5470 => x"94",     5471 => x"93", 
    5472 => x"92",     5473 => x"91",     5474 => x"90",     5475 => x"8E",     5476 => x"8D",     5477 => x"8B",     5478 => x"89",     5479 => x"87", 
    5480 => x"85",     5481 => x"83",     5482 => x"81",     5483 => x"7F",     5484 => x"7D",     5485 => x"7C",     5486 => x"7A",     5487 => x"7A", 
    5488 => x"7A",     5489 => x"7A",     5490 => x"7A",     5491 => x"7A",     5492 => x"7B",     5493 => x"7D",     5494 => x"7F",     5495 => x"80", 
    5496 => x"82",     5497 => x"83",     5498 => x"84",     5499 => x"84",     5500 => x"84",     5501 => x"84",     5502 => x"83",     5503 => x"82", 
    5504 => x"80",     5505 => x"7F",     5506 => x"7E",     5507 => x"7C",     5508 => x"7B",     5509 => x"7B",     5510 => x"7A",     5511 => x"7A", 
    5512 => x"7B",     5513 => x"7C",     5514 => x"7D",     5515 => x"7F",     5516 => x"7F",     5517 => x"80",     5518 => x"82",     5519 => x"84", 
    5520 => x"86",     5521 => x"87",     5522 => x"88",     5523 => x"8A",     5524 => x"8A",     5525 => x"8A",     5526 => x"8B",     5527 => x"8B", 
    5528 => x"8B",     5529 => x"8B",     5530 => x"8B",     5531 => x"8B",     5532 => x"8B",     5533 => x"8A",     5534 => x"8A",     5535 => x"89", 
    5536 => x"89",     5537 => x"89",     5538 => x"89",     5539 => x"8A",     5540 => x"8B",     5541 => x"8C",     5542 => x"8D",     5543 => x"8D", 
    5544 => x"8F",     5545 => x"90",     5546 => x"91",     5547 => x"92",     5548 => x"93",     5549 => x"94",     5550 => x"95",     5551 => x"95", 
    5552 => x"96",     5553 => x"96",     5554 => x"97",     5555 => x"96",     5556 => x"96",     5557 => x"96",     5558 => x"95",     5559 => x"95", 
    5560 => x"94",     5561 => x"92",     5562 => x"91",     5563 => x"8F",     5564 => x"8E",     5565 => x"8C",     5566 => x"8B",     5567 => x"8A", 
    5568 => x"89",     5569 => x"88",     5570 => x"88",     5571 => x"88",     5572 => x"88",     5573 => x"88",     5574 => x"89",     5575 => x"8B", 
    5576 => x"8C",     5577 => x"8E",     5578 => x"8E",     5579 => x"8F",     5580 => x"90",     5581 => x"90",     5582 => x"90",     5583 => x"90", 
    5584 => x"90",     5585 => x"8F",     5586 => x"8F",     5587 => x"8E",     5588 => x"8C",     5589 => x"8B",     5590 => x"8B",     5591 => x"8A", 
    5592 => x"8A",     5593 => x"8A",     5594 => x"8A",     5595 => x"8B",     5596 => x"8B",     5597 => x"8B",     5598 => x"8C",     5599 => x"8C", 
    5600 => x"8C",     5601 => x"8C",     5602 => x"8B",     5603 => x"8B",     5604 => x"8B",     5605 => x"8B",     5606 => x"8A",     5607 => x"8A", 
    5608 => x"89",     5609 => x"88",     5610 => x"87",     5611 => x"86",     5612 => x"86",     5613 => x"86",     5614 => x"86",     5615 => x"86", 
    5616 => x"86",     5617 => x"86",     5618 => x"86",     5619 => x"87",     5620 => x"87",     5621 => x"88",     5622 => x"89",     5623 => x"8A", 
    5624 => x"8B",     5625 => x"8C",     5626 => x"8B",     5627 => x"8A",     5628 => x"89",     5629 => x"88",     5630 => x"88",     5631 => x"87", 
    5632 => x"86",     5633 => x"86",     5634 => x"86",     5635 => x"85",     5636 => x"84",     5637 => x"84",     5638 => x"84",     5639 => x"85", 
    5640 => x"84",     5641 => x"85",     5642 => x"85",     5643 => x"86",     5644 => x"86",     5645 => x"85",     5646 => x"85",     5647 => x"84", 
    5648 => x"84",     5649 => x"83",     5650 => x"83",     5651 => x"82",     5652 => x"80",     5653 => x"7F",     5654 => x"7E",     5655 => x"7D", 
    5656 => x"7C",     5657 => x"7B",     5658 => x"7A",     5659 => x"7A",     5660 => x"7A",     5661 => x"7A",     5662 => x"7B",     5663 => x"7B", 
    5664 => x"7C",     5665 => x"7D",     5666 => x"7D",     5667 => x"7E",     5668 => x"7F",     5669 => x"80",     5670 => x"81",     5671 => x"82", 
    5672 => x"84",     5673 => x"85",     5674 => x"86",     5675 => x"87",     5676 => x"88",     5677 => x"8A",     5678 => x"8B",     5679 => x"8C", 
    5680 => x"8E",     5681 => x"8F",     5682 => x"8F",     5683 => x"90",     5684 => x"90",     5685 => x"90",     5686 => x"90",     5687 => x"90", 
    5688 => x"90",     5689 => x"8F",     5690 => x"8F",     5691 => x"8F",     5692 => x"8F",     5693 => x"90",     5694 => x"90",     5695 => x"90", 
    5696 => x"90",     5697 => x"90",     5698 => x"91",     5699 => x"92",     5700 => x"93",     5701 => x"94",     5702 => x"95",     5703 => x"96", 
    5704 => x"97",     5705 => x"98",     5706 => x"98",     5707 => x"99",     5708 => x"9A",     5709 => x"9B",     5710 => x"9B",     5711 => x"9C", 
    5712 => x"9C",     5713 => x"9B",     5714 => x"9A",     5715 => x"99",     5716 => x"98",     5717 => x"97",     5718 => x"97",     5719 => x"96", 
    5720 => x"95",     5721 => x"94",     5722 => x"92",     5723 => x"91",     5724 => x"90",     5725 => x"8F",     5726 => x"8E",     5727 => x"8E", 
    5728 => x"8E",     5729 => x"8D",     5730 => x"8C",     5731 => x"8C",     5732 => x"8B",     5733 => x"89",     5734 => x"89",     5735 => x"87", 
    5736 => x"86",     5737 => x"86",     5738 => x"85",     5739 => x"84",     5740 => x"83",     5741 => x"83",     5742 => x"83",     5743 => x"82", 
    5744 => x"82",     5745 => x"81",     5746 => x"81",     5747 => x"80",     5748 => x"80",     5749 => x"7F",     5750 => x"7E",     5751 => x"7D", 
    5752 => x"7C",     5753 => x"7B",     5754 => x"7A",     5755 => x"7A",     5756 => x"79",     5757 => x"79",     5758 => x"79",     5759 => x"79", 
    5760 => x"79",     5761 => x"78",     5762 => x"79",     5763 => x"79",     5764 => x"7A",     5765 => x"7B",     5766 => x"7B",     5767 => x"7C", 
    5768 => x"7D",     5769 => x"7F",     5770 => x"80",     5771 => x"81",     5772 => x"82",     5773 => x"83",     5774 => x"84",     5775 => x"86", 
    5776 => x"87",     5777 => x"87",     5778 => x"88",     5779 => x"88",     5780 => x"89",     5781 => x"89",     5782 => x"89",     5783 => x"8A", 
    5784 => x"8A",     5785 => x"8A",     5786 => x"8A",     5787 => x"8A",     5788 => x"8B",     5789 => x"8B",     5790 => x"8B",     5791 => x"8B", 
    5792 => x"8B",     5793 => x"8C",     5794 => x"8D",     5795 => x"8D",     5796 => x"8D",     5797 => x"8E",     5798 => x"8E",     5799 => x"8E", 
    5800 => x"8E",     5801 => x"8E",     5802 => x"8E",     5803 => x"8E",     5804 => x"8E",     5805 => x"8F",     5806 => x"8F",     5807 => x"90", 
    5808 => x"8F",     5809 => x"90",     5810 => x"90",     5811 => x"90",     5812 => x"91",     5813 => x"91",     5814 => x"91",     5815 => x"90", 
    5816 => x"90",     5817 => x"91",     5818 => x"90",     5819 => x"8F",     5820 => x"8E",     5821 => x"8E",     5822 => x"8E",     5823 => x"8E", 
    5824 => x"8F",     5825 => x"8E",     5826 => x"8F",     5827 => x"8F",     5828 => x"8E",     5829 => x"8F",     5830 => x"8F",     5831 => x"8E", 
    5832 => x"8D",     5833 => x"8D",     5834 => x"8E",     5835 => x"8E",     5836 => x"8F",     5837 => x"8F",     5838 => x"8F",     5839 => x"8F", 
    5840 => x"8F",     5841 => x"90",     5842 => x"90",     5843 => x"90",     5844 => x"90",     5845 => x"8F",     5846 => x"8F",     5847 => x"8F", 
    5848 => x"8E",     5849 => x"8E",     5850 => x"8C",     5851 => x"8C",     5852 => x"8B",     5853 => x"8B",     5854 => x"8A",     5855 => x"89", 
    5856 => x"88",     5857 => x"88",     5858 => x"88",     5859 => x"88",     5860 => x"88",     5861 => x"87",     5862 => x"86",     5863 => x"86", 
    5864 => x"87",     5865 => x"88",     5866 => x"88",     5867 => x"88",     5868 => x"87",     5869 => x"87",     5870 => x"87",     5871 => x"87", 
    5872 => x"86",     5873 => x"86",     5874 => x"85",     5875 => x"84",     5876 => x"84",     5877 => x"83",     5878 => x"82",     5879 => x"81", 
    5880 => x"80",     5881 => x"7F",     5882 => x"7F",     5883 => x"7F",     5884 => x"7F",     5885 => x"7F",     5886 => x"7E",     5887 => x"7E", 
    5888 => x"7E",     5889 => x"7E",     5890 => x"7F",     5891 => x"80",     5892 => x"81",     5893 => x"81",     5894 => x"82",     5895 => x"83", 
    5896 => x"83",     5897 => x"83",     5898 => x"82",     5899 => x"82",     5900 => x"83",     5901 => x"83",     5902 => x"83",     5903 => x"83", 
    5904 => x"82",     5905 => x"82",     5906 => x"81",     5907 => x"81",     5908 => x"81",     5909 => x"81",     5910 => x"80",     5911 => x"80", 
    5912 => x"7F",     5913 => x"7F",     5914 => x"7E",     5915 => x"7D",     5916 => x"7D",     5917 => x"7E",     5918 => x"7E",     5919 => x"7F", 
    5920 => x"7F",     5921 => x"7F",     5922 => x"80",     5923 => x"81",     5924 => x"82",     5925 => x"83",     5926 => x"83",     5927 => x"84", 
    5928 => x"85",     5929 => x"86",     5930 => x"87",     5931 => x"88",     5932 => x"89",     5933 => x"8A",     5934 => x"8B",     5935 => x"8C", 
    5936 => x"8D",     5937 => x"8D",     5938 => x"8D",     5939 => x"8E",     5940 => x"8E",     5941 => x"8F",     5942 => x"90",     5943 => x"90", 
    5944 => x"91",     5945 => x"92",     5946 => x"92",     5947 => x"93",     5948 => x"94",     5949 => x"95",     5950 => x"97",     5951 => x"97", 
    5952 => x"98",     5953 => x"98",     5954 => x"99",     5955 => x"9A",     5956 => x"9A",     5957 => x"9A",     5958 => x"9A",     5959 => x"9B", 
    5960 => x"9C",     5961 => x"9D",     5962 => x"9D",     5963 => x"9D",     5964 => x"9D",     5965 => x"9C",     5966 => x"9B",     5967 => x"9A", 
    5968 => x"99",     5969 => x"99",     5970 => x"97",     5971 => x"97",     5972 => x"96",     5973 => x"95",     5974 => x"94",     5975 => x"93", 
    5976 => x"93",     5977 => x"92",     5978 => x"92",     5979 => x"92",     5980 => x"92",     5981 => x"93",     5982 => x"93",     5983 => x"92", 
    5984 => x"92",     5985 => x"91",     5986 => x"91",     5987 => x"90",     5988 => x"90",     5989 => x"90",     5990 => x"8F",     5991 => x"8E", 
    5992 => x"8D",     5993 => x"8C",     5994 => x"8B",     5995 => x"8A",     5996 => x"8A",     5997 => x"89",     5998 => x"89",     5999 => x"88", 
    6000 => x"88",     6001 => x"88",     6002 => x"87",     6003 => x"87",     6004 => x"86",     6005 => x"86",     6006 => x"85",     6007 => x"85", 
    6008 => x"85",     6009 => x"84",     6010 => x"84",     6011 => x"84",     6012 => x"84",     6013 => x"83",     6014 => x"82",     6015 => x"82", 
    6016 => x"81",     6017 => x"81",     6018 => x"81",     6019 => x"81",     6020 => x"81",     6021 => x"80",     6022 => x"7F",     6023 => x"7F", 
    6024 => x"7E",     6025 => x"7D",     6026 => x"7C",     6027 => x"7C",     6028 => x"7B",     6029 => x"7B",     6030 => x"7A",     6031 => x"7A", 
    6032 => x"78",     6033 => x"78",     6034 => x"77",     6035 => x"78",     6036 => x"78",     6037 => x"79",     6038 => x"79",     6039 => x"7A", 
    6040 => x"7C",     6041 => x"7D",     6042 => x"7E",     6043 => x"7F",     6044 => x"7F",     6045 => x"80",     6046 => x"80",     6047 => x"81", 
    6048 => x"81",     6049 => x"81",     6050 => x"81",     6051 => x"80",     6052 => x"80",     6053 => x"80",     6054 => x"7F",     6055 => x"7E", 
    6056 => x"7E",     6057 => x"7F",     6058 => x"7F",     6059 => x"7F",     6060 => x"80",     6061 => x"81",     6062 => x"82",     6063 => x"83", 
    6064 => x"83",     6065 => x"85",     6066 => x"86",     6067 => x"87",     6068 => x"87",     6069 => x"88",     6070 => x"89",     6071 => x"89", 
    6072 => x"8A",     6073 => x"8A",     6074 => x"8A",     6075 => x"8A",     6076 => x"8A",     6077 => x"8A",     6078 => x"8B",     6079 => x"8C", 
    6080 => x"8C",     6081 => x"8D",     6082 => x"8E",     6083 => x"8E",     6084 => x"8F",     6085 => x"90",     6086 => x"91",     6087 => x"92", 
    6088 => x"92",     6089 => x"93",     6090 => x"94",     6091 => x"94",     6092 => x"95",     6093 => x"94",     6094 => x"94",     6095 => x"95", 
    6096 => x"95",     6097 => x"96",     6098 => x"97",     6099 => x"97",     6100 => x"98",     6101 => x"99",     6102 => x"9A",     6103 => x"9B", 
    6104 => x"9C",     6105 => x"9C",     6106 => x"9D",     6107 => x"9D",     6108 => x"9D",     6109 => x"9D",     6110 => x"9D",     6111 => x"9C", 
    6112 => x"9C",     6113 => x"9B",     6114 => x"9A",     6115 => x"99",     6116 => x"97",     6117 => x"96",     6118 => x"94",     6119 => x"93", 
    6120 => x"92",     6121 => x"91",     6122 => x"90",     6123 => x"8F",     6124 => x"8E",     6125 => x"8E",     6126 => x"8D",     6127 => x"8C", 
    6128 => x"8C",     6129 => x"8C",     6130 => x"8C",     6131 => x"8B",     6132 => x"8B",     6133 => x"8B",     6134 => x"8B",     6135 => x"8B", 
    6136 => x"8B",     6137 => x"8B",     6138 => x"8A",     6139 => x"8A",     6140 => x"8A",     6141 => x"89",     6142 => x"89",     6143 => x"88", 
    6144 => x"87",     6145 => x"86",     6146 => x"86",     6147 => x"85",     6148 => x"85",     6149 => x"84",     6150 => x"83",     6151 => x"82", 
    6152 => x"81",     6153 => x"80",     6154 => x"80",     6155 => x"7F",     6156 => x"7E",     6157 => x"7D",     6158 => x"7D",     6159 => x"7C", 
    6160 => x"7C",     6161 => x"7C",     6162 => x"7C",     6163 => x"7C",     6164 => x"7C",     6165 => x"7C",     6166 => x"7B",     6167 => x"7B", 
    6168 => x"7B",     6169 => x"7C",     6170 => x"7C",     6171 => x"7C",     6172 => x"7C",     6173 => x"7C",     6174 => x"7C",     6175 => x"7B", 
    6176 => x"7B",     6177 => x"7B",     6178 => x"7B",     6179 => x"7B",     6180 => x"7B",     6181 => x"7B",     6182 => x"7B",     6183 => x"7B", 
    6184 => x"7B",     6185 => x"7C",     6186 => x"7C",     6187 => x"7D",     6188 => x"7E",     6189 => x"7E",     6190 => x"7F",     6191 => x"80", 
    6192 => x"81",     6193 => x"82",     6194 => x"84",     6195 => x"85",     6196 => x"86",     6197 => x"87",     6198 => x"89",     6199 => x"8A", 
    6200 => x"8C",     6201 => x"8D",     6202 => x"8E",     6203 => x"8F",     6204 => x"90",     6205 => x"90",     6206 => x"91",     6207 => x"91", 
    6208 => x"92",     6209 => x"92",     6210 => x"93",     6211 => x"93",     6212 => x"93",     6213 => x"93",     6214 => x"92",     6215 => x"92", 
    6216 => x"92",     6217 => x"91",     6218 => x"91",     6219 => x"91",     6220 => x"91",     6221 => x"91",     6222 => x"91",     6223 => x"91", 
    6224 => x"90",     6225 => x"91",     6226 => x"92",     6227 => x"93",     6228 => x"93",     6229 => x"94",     6230 => x"94",     6231 => x"95", 
    6232 => x"95",     6233 => x"95",     6234 => x"96",     6235 => x"97",     6236 => x"97",     6237 => x"97",     6238 => x"97",     6239 => x"97", 
    6240 => x"96",     6241 => x"96",     6242 => x"95",     6243 => x"95",     6244 => x"95",     6245 => x"94",     6246 => x"94",     6247 => x"93", 
    6248 => x"92",     6249 => x"92",     6250 => x"91",     6251 => x"90",     6252 => x"8F",     6253 => x"8E",     6254 => x"8E",     6255 => x"8E", 
    6256 => x"8D",     6257 => x"8C",     6258 => x"8B",     6259 => x"8B",     6260 => x"8A",     6261 => x"89",     6262 => x"88",     6263 => x"88", 
    6264 => x"88",     6265 => x"87",     6266 => x"87",     6267 => x"86",     6268 => x"84",     6269 => x"83",     6270 => x"83",     6271 => x"82", 
    6272 => x"82",     6273 => x"82",     6274 => x"82",     6275 => x"81",     6276 => x"80",     6277 => x"80",     6278 => x"7F",     6279 => x"7F", 
    6280 => x"7F",     6281 => x"7F",     6282 => x"7F",     6283 => x"80",     6284 => x"80",     6285 => x"7F",     6286 => x"7F",     6287 => x"7F", 
    6288 => x"80",     6289 => x"80",     6290 => x"80",     6291 => x"81",     6292 => x"81",     6293 => x"81",     6294 => x"81",     6295 => x"82", 
    6296 => x"82",     6297 => x"82",     6298 => x"82",     6299 => x"83",     6300 => x"83",     6301 => x"83",     6302 => x"83",     6303 => x"84", 
    6304 => x"84",     6305 => x"84",     6306 => x"84",     6307 => x"84",     6308 => x"84",     6309 => x"84",     6310 => x"84",     6311 => x"84", 
    6312 => x"84",     6313 => x"85",     6314 => x"85",     6315 => x"85",     6316 => x"85",     6317 => x"85",     6318 => x"85",     6319 => x"85", 
    6320 => x"86",     6321 => x"86",     6322 => x"87",     6323 => x"88",     6324 => x"88",     6325 => x"89",     6326 => x"8A",     6327 => x"8A", 
    6328 => x"8A",     6329 => x"8A",     6330 => x"8B",     6331 => x"8C",     6332 => x"8C",     6333 => x"8C",     6334 => x"8D",     6335 => x"8D", 
    6336 => x"8D",     6337 => x"8E",     6338 => x"8E",     6339 => x"8E",     6340 => x"8E",     6341 => x"8E",     6342 => x"8E",     6343 => x"8F", 
    6344 => x"8F",     6345 => x"8F",     6346 => x"8F",     6347 => x"8F",     6348 => x"8E",     6349 => x"8E",     6350 => x"8D",     6351 => x"8D", 
    6352 => x"8D",     6353 => x"8C",     6354 => x"8C",     6355 => x"8C",     6356 => x"8D",     6357 => x"8C",     6358 => x"8C",     6359 => x"8C", 
    6360 => x"8C",     6361 => x"8C",     6362 => x"8C",     6363 => x"8C",     6364 => x"8C",     6365 => x"8C",     6366 => x"8C",     6367 => x"8C", 
    6368 => x"8C",     6369 => x"8C",     6370 => x"8C",     6371 => x"8B",     6372 => x"8B",     6373 => x"8B",     6374 => x"8B",     6375 => x"8A", 
    6376 => x"8A",     6377 => x"8A",     6378 => x"89",     6379 => x"89",     6380 => x"89",     6381 => x"88",     6382 => x"88",     6383 => x"88", 
    6384 => x"87",     6385 => x"87",     6386 => x"87",     6387 => x"87",     6388 => x"87",     6389 => x"87",     6390 => x"87",     6391 => x"87", 
    6392 => x"87",     6393 => x"88",     6394 => x"89",     6395 => x"89",     6396 => x"8A",     6397 => x"8B",     6398 => x"8B",     6399 => x"8C", 
    6400 => x"8D",     6401 => x"8D",     6402 => x"8E",     6403 => x"8E",     6404 => x"8F",     6405 => x"8E",     6406 => x"8E",     6407 => x"8E", 
    6408 => x"8E",     6409 => x"8E",     6410 => x"8E",     6411 => x"8D",     6412 => x"8D",     6413 => x"8C",     6414 => x"8B",     6415 => x"8B", 
    6416 => x"8A",     6417 => x"8A",     6418 => x"8A",     6419 => x"8A",     6420 => x"8A",     6421 => x"8A",     6422 => x"8A",     6423 => x"8A", 
    6424 => x"8A",     6425 => x"8B",     6426 => x"8C",     6427 => x"8C",     6428 => x"8C",     6429 => x"8D",     6430 => x"8C",     6431 => x"8C", 
    6432 => x"8C",     6433 => x"8B",     6434 => x"8B",     6435 => x"8B",     6436 => x"8B",     6437 => x"8A",     6438 => x"89",     6439 => x"89", 
    6440 => x"88",     6441 => x"87",     6442 => x"87",     6443 => x"86",     6444 => x"86",     6445 => x"85",     6446 => x"85",     6447 => x"85", 
    6448 => x"84",     6449 => x"84",     6450 => x"84",     6451 => x"84",     6452 => x"84",     6453 => x"84",     6454 => x"85",     6455 => x"85", 
    6456 => x"85",     6457 => x"85",     6458 => x"85",     6459 => x"85",     6460 => x"84",     6461 => x"85",     6462 => x"85",     6463 => x"86", 
    6464 => x"85",     6465 => x"85",     6466 => x"84",     6467 => x"83",     6468 => x"83",     6469 => x"82",     6470 => x"82",     6471 => x"82", 
    6472 => x"82",     6473 => x"81",     6474 => x"80",     6475 => x"80",     6476 => x"7F",     6477 => x"7F",     6478 => x"7F",     6479 => x"80", 
    6480 => x"81",     6481 => x"81",     6482 => x"82",     6483 => x"83",     6484 => x"83",     6485 => x"84",     6486 => x"84",     6487 => x"84", 
    6488 => x"85",     6489 => x"86",     6490 => x"87",     6491 => x"88",     6492 => x"89",     6493 => x"8A",     6494 => x"8A",     6495 => x"8B", 
    6496 => x"8B",     6497 => x"8C",     6498 => x"8D",     6499 => x"8E",     6500 => x"8E",     6501 => x"8F",     6502 => x"8F",     6503 => x"90", 
    6504 => x"90",     6505 => x"90",     6506 => x"91",     6507 => x"91",     6508 => x"91",     6509 => x"92",     6510 => x"92",     6511 => x"92", 
    6512 => x"92",     6513 => x"92",     6514 => x"92",     6515 => x"92",     6516 => x"92",     6517 => x"93",     6518 => x"93",     6519 => x"93", 
    6520 => x"93",     6521 => x"93",     6522 => x"94",     6523 => x"94",     6524 => x"94",     6525 => x"94",     6526 => x"94",     6527 => x"95", 
    6528 => x"95",     6529 => x"95",     6530 => x"95",     6531 => x"96",     6532 => x"96",     6533 => x"96",     6534 => x"96",     6535 => x"97", 
    6536 => x"97",     6537 => x"97",     6538 => x"96",     6539 => x"94",     6540 => x"93",     6541 => x"93",     6542 => x"91",     6543 => x"90", 
    6544 => x"8F",     6545 => x"8E",     6546 => x"8D",     6547 => x"8C",     6548 => x"8A",     6549 => x"89",     6550 => x"88",     6551 => x"87", 
    6552 => x"85",     6553 => x"84",     6554 => x"84",     6555 => x"83",     6556 => x"82",     6557 => x"81",     6558 => x"80",     6559 => x"80", 
    6560 => x"80",     6561 => x"80",     6562 => x"80",     6563 => x"81",     6564 => x"81",     6565 => x"81",     6566 => x"82",     6567 => x"82", 
    6568 => x"82",     6569 => x"83",     6570 => x"83",     6571 => x"83",     6572 => x"83",     6573 => x"83",     6574 => x"83",     6575 => x"83", 
    6576 => x"82",     6577 => x"82",     6578 => x"82",     6579 => x"82",     6580 => x"81",     6581 => x"80",     6582 => x"7F",     6583 => x"7E", 
    6584 => x"7E",     6585 => x"7D",     6586 => x"7C",     6587 => x"7C",     6588 => x"7C",     6589 => x"7B",     6590 => x"7B",     6591 => x"7A", 
    6592 => x"7A",     6593 => x"7A",     6594 => x"7A",     6595 => x"7A",     6596 => x"7A",     6597 => x"7B",     6598 => x"7C",     6599 => x"7C", 
    6600 => x"7C",     6601 => x"7C",     6602 => x"7C",     6603 => x"7C",     6604 => x"7C",     6605 => x"7D",     6606 => x"7E",     6607 => x"7F", 
    6608 => x"80",     6609 => x"80",     6610 => x"81",     6611 => x"81",     6612 => x"82",     6613 => x"82",     6614 => x"83",     6615 => x"84", 
    6616 => x"85",     6617 => x"86",     6618 => x"87",     6619 => x"88",     6620 => x"89",     6621 => x"8B",     6622 => x"8C",     6623 => x"8D", 
    6624 => x"8D",     6625 => x"8E",     6626 => x"8E",     6627 => x"8F",     6628 => x"90",     6629 => x"91",     6630 => x"91",     6631 => x"92", 
    6632 => x"92",     6633 => x"92",     6634 => x"92",     6635 => x"93",     6636 => x"93",     6637 => x"94",     6638 => x"95",     6639 => x"96", 
    6640 => x"97",     6641 => x"98",     6642 => x"98",     6643 => x"99",     6644 => x"9A",     6645 => x"9A",     6646 => x"9B",     6647 => x"9C", 
    6648 => x"9C",     6649 => x"9D",     6650 => x"9E",     6651 => x"9E",     6652 => x"9E",     6653 => x"9E",     6654 => x"9E",     6655 => x"9D", 
    6656 => x"9D",     6657 => x"9C",     6658 => x"9C",     6659 => x"9B",     6660 => x"9A",     6661 => x"99",     6662 => x"98",     6663 => x"98", 
    6664 => x"98",     6665 => x"96",     6666 => x"95",     6667 => x"94",     6668 => x"93",     6669 => x"92",     6670 => x"91",     6671 => x"90", 
    6672 => x"90",     6673 => x"8F",     6674 => x"8E",     6675 => x"8D",     6676 => x"8C",     6677 => x"8B",     6678 => x"8A",     6679 => x"8A", 
    6680 => x"8A",     6681 => x"89",     6682 => x"89",     6683 => x"88",     6684 => x"88",     6685 => x"87",     6686 => x"87",     6687 => x"86", 
    6688 => x"86",     6689 => x"86",     6690 => x"85",     6691 => x"85",     6692 => x"84",     6693 => x"84",     6694 => x"83",     6695 => x"82", 
    6696 => x"81",     6697 => x"81",     6698 => x"80",     6699 => x"80",     6700 => x"80",     6701 => x"80",     6702 => x"7F",     6703 => x"7F", 
    6704 => x"7E",     6705 => x"7E",     6706 => x"7D",     6707 => x"7C",     6708 => x"7C",     6709 => x"7C",     6710 => x"7C",     6711 => x"7C", 
    6712 => x"7C",     6713 => x"7C",     6714 => x"7B",     6715 => x"7B",     6716 => x"7A",     6717 => x"7A",     6718 => x"7A",     6719 => x"7A", 
    6720 => x"7B",     6721 => x"7B",     6722 => x"7C",     6723 => x"7C",     6724 => x"7D",     6725 => x"7D",     6726 => x"7D",     6727 => x"7E", 
    6728 => x"7F",     6729 => x"7F",     6730 => x"80",     6731 => x"80",     6732 => x"80",     6733 => x"80",     6734 => x"80",     6735 => x"80", 
    6736 => x"81",     6737 => x"81",     6738 => x"82",     6739 => x"82",     6740 => x"83",     6741 => x"83",     6742 => x"84",     6743 => x"84", 
    6744 => x"85",     6745 => x"85",     6746 => x"86",     6747 => x"87",     6748 => x"87",     6749 => x"87",     6750 => x"87",     6751 => x"87", 
    6752 => x"87",     6753 => x"87",     6754 => x"86",     6755 => x"87",     6756 => x"87",     6757 => x"87",     6758 => x"87",     6759 => x"87", 
    6760 => x"88",     6761 => x"88",     6762 => x"88",     6763 => x"89",     6764 => x"89",     6765 => x"8A",     6766 => x"8B",     6767 => x"8D", 
    6768 => x"8E",     6769 => x"8E",     6770 => x"8F",     6771 => x"8F",     6772 => x"90",     6773 => x"90",     6774 => x"91",     6775 => x"92", 
    6776 => x"92",     6777 => x"93",     6778 => x"93",     6779 => x"93",     6780 => x"94",     6781 => x"94",     6782 => x"94",     6783 => x"94", 
    6784 => x"93",     6785 => x"93",     6786 => x"93",     6787 => x"94",     6788 => x"94",     6789 => x"93",     6790 => x"93",     6791 => x"93", 
    6792 => x"93",     6793 => x"93",     6794 => x"93",     6795 => x"93",     6796 => x"93",     6797 => x"93",     6798 => x"92",     6799 => x"92", 
    6800 => x"91",     6801 => x"91",     6802 => x"91",     6803 => x"90",     6804 => x"90",     6805 => x"90",     6806 => x"90",     6807 => x"90", 
    6808 => x"90",     6809 => x"90",     6810 => x"90",     6811 => x"90",     6812 => x"8F",     6813 => x"8F",     6814 => x"8F",     6815 => x"8F", 
    6816 => x"8E",     6817 => x"8E",     6818 => x"8D",     6819 => x"8D",     6820 => x"8C",     6821 => x"8C",     6822 => x"8C",     6823 => x"8B", 
    6824 => x"8B",     6825 => x"8B",     6826 => x"8B",     6827 => x"8B",     6828 => x"8C",     6829 => x"8C",     6830 => x"8C",     6831 => x"8B", 
    6832 => x"8B",     6833 => x"8A",     6834 => x"8A",     6835 => x"89",     6836 => x"89",     6837 => x"89",     6838 => x"88",     6839 => x"88", 
    6840 => x"87",     6841 => x"86",     6842 => x"84",     6843 => x"83",     6844 => x"82",     6845 => x"82",     6846 => x"82",     6847 => x"82", 
    6848 => x"82",     6849 => x"81",     6850 => x"80",     6851 => x"7F",     6852 => x"7E",     6853 => x"7E",     6854 => x"7E",     6855 => x"7E", 
    6856 => x"7F",     6857 => x"7F",     6858 => x"7F",     6859 => x"7F",     6860 => x"80",     6861 => x"7F",     6862 => x"7F",     6863 => x"7F", 
    6864 => x"80",     6865 => x"80",     6866 => x"80",     6867 => x"80",     6868 => x"80",     6869 => x"80",     6870 => x"80",     6871 => x"80", 
    6872 => x"7F",     6873 => x"7F",     6874 => x"7F",     6875 => x"7F",     6876 => x"7F",     6877 => x"7F",     6878 => x"7F",     6879 => x"7E", 
    6880 => x"7E",     6881 => x"7E",     6882 => x"7E",     6883 => x"7F",     6884 => x"80",     6885 => x"81",     6886 => x"82",     6887 => x"83", 
    6888 => x"83",     6889 => x"84",     6890 => x"85",     6891 => x"86",     6892 => x"88",     6893 => x"89",     6894 => x"8A",     6895 => x"8A", 
    6896 => x"8A",     6897 => x"8A",     6898 => x"8B",     6899 => x"8B",     6900 => x"8C",     6901 => x"8C",     6902 => x"8D",     6903 => x"8F", 
    6904 => x"90",     6905 => x"91",     6906 => x"91",     6907 => x"91",     6908 => x"92",     6909 => x"92",     6910 => x"93",     6911 => x"94", 
    6912 => x"94",     6913 => x"95",     6914 => x"96",     6915 => x"96",     6916 => x"96",     6917 => x"96",     6918 => x"96",     6919 => x"96", 
    6920 => x"95",     6921 => x"95",     6922 => x"95",     6923 => x"95",     6924 => x"96",     6925 => x"96",     6926 => x"96",     6927 => x"96", 
    6928 => x"96",     6929 => x"96",     6930 => x"96",     6931 => x"96",     6932 => x"97",     6933 => x"96",     6934 => x"97",     6935 => x"97", 
    6936 => x"97",     6937 => x"96",     6938 => x"96",     6939 => x"95",     6940 => x"94",     6941 => x"94",     6942 => x"93",     6943 => x"93", 
    6944 => x"92",     6945 => x"92",     6946 => x"91",     6947 => x"90",     6948 => x"8F",     6949 => x"8F",     6950 => x"8E",     6951 => x"8E", 
    6952 => x"8E",     6953 => x"8E",     6954 => x"8D",     6955 => x"8D",     6956 => x"8D",     6957 => x"8D",     6958 => x"8C",     6959 => x"8B", 
    6960 => x"8A",     6961 => x"89",     6962 => x"88",     6963 => x"88",     6964 => x"87",     6965 => x"87",     6966 => x"86",     6967 => x"85", 
    6968 => x"84",     6969 => x"84",     6970 => x"83",     6971 => x"83",     6972 => x"83",     6973 => x"83",     6974 => x"83",     6975 => x"82", 
    6976 => x"81",     6977 => x"80",     6978 => x"7F",     6979 => x"7F",     6980 => x"7E",     6981 => x"7F",     6982 => x"7F",     6983 => x"7E", 
    6984 => x"7E",     6985 => x"7D",     6986 => x"7C",     6987 => x"7B",     6988 => x"7B",     6989 => x"7A",     6990 => x"7A",     6991 => x"7A", 
    6992 => x"7B",     6993 => x"7B",     6994 => x"7B",     6995 => x"7B",     6996 => x"7B",     6997 => x"7B",     6998 => x"7B",     6999 => x"7C", 
    7000 => x"7C",     7001 => x"7D",     7002 => x"7D",     7003 => x"7D",     7004 => x"7D",     7005 => x"7D",     7006 => x"7D",     7007 => x"7D", 
    7008 => x"7D",     7009 => x"7E",     7010 => x"7E",     7011 => x"7F",     7012 => x"7F",     7013 => x"7F",     7014 => x"80",     7015 => x"80", 
    7016 => x"81",     7017 => x"81",     7018 => x"82",     7019 => x"82",     7020 => x"83",     7021 => x"83",     7022 => x"84",     7023 => x"84", 
    7024 => x"85",     7025 => x"85",     7026 => x"87",     7027 => x"88",     7028 => x"8A",     7029 => x"8B",     7030 => x"8D",     7031 => x"8E", 
    7032 => x"8F",     7033 => x"90",     7034 => x"91",     7035 => x"92",     7036 => x"93",     7037 => x"94",     7038 => x"94",     7039 => x"95", 
    7040 => x"96",     7041 => x"96",     7042 => x"96",     7043 => x"96",     7044 => x"95",     7045 => x"96",     7046 => x"96",     7047 => x"96", 
    7048 => x"97",     7049 => x"97",     7050 => x"96",     7051 => x"96",     7052 => x"95",     7053 => x"95",     7054 => x"95",     7055 => x"94", 
    7056 => x"94",     7057 => x"95",     7058 => x"95",     7059 => x"95",     7060 => x"95",     7061 => x"95",     7062 => x"95",     7063 => x"95", 
    7064 => x"94",     7065 => x"95",     7066 => x"95",     7067 => x"95",     7068 => x"94",     7069 => x"94",     7070 => x"93",     7071 => x"93", 
    7072 => x"92",     7073 => x"92",     7074 => x"92",     7075 => x"92",     7076 => x"92",     7077 => x"92",     7078 => x"91",     7079 => x"90", 
    7080 => x"8F",     7081 => x"8F",     7082 => x"8F",     7083 => x"8E",     7084 => x"8E",     7085 => x"8D",     7086 => x"8D",     7087 => x"8C", 
    7088 => x"8C",     7089 => x"8B",     7090 => x"8A",     7091 => x"8A",     7092 => x"8A",     7093 => x"8A",     7094 => x"89",     7095 => x"89", 
    7096 => x"89",     7097 => x"89",     7098 => x"88",     7099 => x"88",     7100 => x"87",     7101 => x"86",     7102 => x"86",     7103 => x"86", 
    7104 => x"86",     7105 => x"86",     7106 => x"85",     7107 => x"84",     7108 => x"84",     7109 => x"83",     7110 => x"82",     7111 => x"81", 
    7112 => x"80",     7113 => x"80",     7114 => x"7F",     7115 => x"7E",     7116 => x"7D",     7117 => x"7D",     7118 => x"7C",     7119 => x"7C", 
    7120 => x"7C",     7121 => x"7C",     7122 => x"7C",     7123 => x"7C",     7124 => x"7C",     7125 => x"7C",     7126 => x"7C",     7127 => x"7C", 
    7128 => x"7C",     7129 => x"7C",     7130 => x"7C",     7131 => x"7D",     7132 => x"7D",     7133 => x"7D",     7134 => x"7D",     7135 => x"7D", 
    7136 => x"7D",     7137 => x"7D",     7138 => x"7D",     7139 => x"7D",     7140 => x"7D",     7141 => x"7D",     7142 => x"7E",     7143 => x"7E", 
    7144 => x"7E",     7145 => x"7F",     7146 => x"7F",     7147 => x"80",     7148 => x"80",     7149 => x"80",     7150 => x"80",     7151 => x"80", 
    7152 => x"81",     7153 => x"82",     7154 => x"83",     7155 => x"84",     7156 => x"84",     7157 => x"85",     7158 => x"86",     7159 => x"86", 
    7160 => x"87",     7161 => x"87",     7162 => x"88",     7163 => x"8A",     7164 => x"8B",     7165 => x"8D",     7166 => x"8D",     7167 => x"8E", 
    7168 => x"8E",     7169 => x"8F",     7170 => x"90",     7171 => x"90",     7172 => x"92",     7173 => x"92",     7174 => x"93",     7175 => x"94", 
    7176 => x"95",     7177 => x"95",     7178 => x"95",     7179 => x"95",     7180 => x"96",     7181 => x"96",     7182 => x"97",     7183 => x"97", 
    7184 => x"97",     7185 => x"97",     7186 => x"97",     7187 => x"98",     7188 => x"98",     7189 => x"98",     7190 => x"98",     7191 => x"98", 
    7192 => x"98",     7193 => x"98",     7194 => x"98",     7195 => x"98",     7196 => x"98",     7197 => x"99",     7198 => x"98",     7199 => x"98", 
    7200 => x"98",     7201 => x"98",     7202 => x"98",     7203 => x"98",     7204 => x"98",     7205 => x"98",     7206 => x"98",     7207 => x"97", 
    7208 => x"98",     7209 => x"97",     7210 => x"97",     7211 => x"97",     7212 => x"96",     7213 => x"96",     7214 => x"94",     7215 => x"93", 
    7216 => x"93",     7217 => x"92",     7218 => x"91",     7219 => x"90",     7220 => x"8E",     7221 => x"8D",     7222 => x"8C",     7223 => x"8B", 
    7224 => x"89",     7225 => x"88",     7226 => x"87",     7227 => x"87",     7228 => x"86",     7229 => x"84",     7230 => x"83",     7231 => x"82", 
    7232 => x"81",     7233 => x"80",     7234 => x"7F",     7235 => x"7F",     7236 => x"7F",     7237 => x"7E",     7238 => x"7E",     7239 => x"7D", 
    7240 => x"7D",     7241 => x"7D",     7242 => x"7D",     7243 => x"7C",     7244 => x"7C",     7245 => x"7C",     7246 => x"7C",     7247 => x"7C", 
    7248 => x"7C",     7249 => x"7C",     7250 => x"7C",     7251 => x"7D",     7252 => x"7D",     7253 => x"7D",     7254 => x"7E",     7255 => x"7E", 
    7256 => x"7F",     7257 => x"7F",     7258 => x"7F",     7259 => x"7F",     7260 => x"80",     7261 => x"80",     7262 => x"81",     7263 => x"81", 
    7264 => x"81",     7265 => x"81",     7266 => x"81",     7267 => x"81",     7268 => x"80",     7269 => x"80",     7270 => x"80",     7271 => x"80", 
    7272 => x"7F",     7273 => x"7F",     7274 => x"7F",     7275 => x"7F",     7276 => x"80",     7277 => x"80",     7278 => x"7F",     7279 => x"7F", 
    7280 => x"7E",     7281 => x"7F",     7282 => x"7F",     7283 => x"7E",     7284 => x"7F",     7285 => x"7F",     7286 => x"7F",     7287 => x"80", 
    7288 => x"81",     7289 => x"81",     7290 => x"82",     7291 => x"83",     7292 => x"84",     7293 => x"85",     7294 => x"85",     7295 => x"86", 
    7296 => x"88",     7297 => x"88",     7298 => x"89",     7299 => x"89",     7300 => x"8A",     7301 => x"8A",     7302 => x"8A",     7303 => x"8B", 
    7304 => x"8C",     7305 => x"8C",     7306 => x"8D",     7307 => x"8D",     7308 => x"8D",     7309 => x"8D",     7310 => x"8E",     7311 => x"8E", 
    7312 => x"8E",     7313 => x"8E",     7314 => x"8F",     7315 => x"8F",     7316 => x"90",     7317 => x"91",     7318 => x"91",     7319 => x"92", 
    7320 => x"92",     7321 => x"93",     7322 => x"94",     7323 => x"94",     7324 => x"94",     7325 => x"94",     7326 => x"95",     7327 => x"95", 
    7328 => x"95",     7329 => x"95",     7330 => x"96",     7331 => x"97",     7332 => x"97",     7333 => x"98",     7334 => x"98",     7335 => x"98", 
    7336 => x"98",     7337 => x"99",     7338 => x"99",     7339 => x"9A",     7340 => x"99",     7341 => x"99",     7342 => x"9A",     7343 => x"99", 
    7344 => x"99",     7345 => x"99",     7346 => x"99",     7347 => x"99",     7348 => x"98",     7349 => x"99",     7350 => x"99",     7351 => x"99", 
    7352 => x"97",     7353 => x"97",     7354 => x"96",     7355 => x"96",     7356 => x"95",     7357 => x"94",     7358 => x"93",     7359 => x"92", 
    7360 => x"91",     7361 => x"90",     7362 => x"8F",     7363 => x"8E",     7364 => x"8D",     7365 => x"8C",     7366 => x"8B",     7367 => x"89", 
    7368 => x"88",     7369 => x"87",     7370 => x"86",     7371 => x"85",     7372 => x"85",     7373 => x"83",     7374 => x"83",     7375 => x"83", 
    7376 => x"82",     7377 => x"81",     7378 => x"81",     7379 => x"81",     7380 => x"80",     7381 => x"7F",     7382 => x"7F",     7383 => x"7E", 
    7384 => x"7E",     7385 => x"7E",     7386 => x"7E",     7387 => x"7E",     7388 => x"7D",     7389 => x"7D",     7390 => x"7D",     7391 => x"7C", 
    7392 => x"7B",     7393 => x"7B",     7394 => x"7A",     7395 => x"7A",     7396 => x"7A",     7397 => x"79",     7398 => x"78",     7399 => x"78", 
    7400 => x"78",     7401 => x"78",     7402 => x"78",     7403 => x"77",     7404 => x"77",     7405 => x"76",     7406 => x"77",     7407 => x"76", 
    7408 => x"76",     7409 => x"76",     7410 => x"76",     7411 => x"77",     7412 => x"77",     7413 => x"76",     7414 => x"77",     7415 => x"78", 
    7416 => x"79",     7417 => x"79",     7418 => x"7A",     7419 => x"7A",     7420 => x"7B",     7421 => x"7C",     7422 => x"7D",     7423 => x"7D", 
    7424 => x"7E",     7425 => x"7F",     7426 => x"81",     7427 => x"82",     7428 => x"82",     7429 => x"82",     7430 => x"84",     7431 => x"85", 
    7432 => x"86",     7433 => x"87",     7434 => x"87",     7435 => x"88",     7436 => x"8A",     7437 => x"8A",     7438 => x"8A",     7439 => x"8A", 
    7440 => x"8C",     7441 => x"8E",     7442 => x"8E",     7443 => x"90",     7444 => x"90",     7445 => x"91",     7446 => x"92",     7447 => x"93", 
    7448 => x"94",     7449 => x"95",     7450 => x"96",     7451 => x"97",     7452 => x"97",     7453 => x"99",     7454 => x"9B",     7455 => x"9C", 
    7456 => x"9C",     7457 => x"9B",     7458 => x"9C",     7459 => x"9D",     7460 => x"9D",     7461 => x"9D",     7462 => x"9D",     7463 => x"9D", 
    7464 => x"9D",     7465 => x"9D",     7466 => x"9C",     7467 => x"9C",     7468 => x"9C",     7469 => x"9A",     7470 => x"9A",     7471 => x"9A", 
    7472 => x"99",     7473 => x"99",     7474 => x"99",     7475 => x"98",     7476 => x"98",     7477 => x"97",     7478 => x"97",     7479 => x"97", 
    7480 => x"96",     7481 => x"95",     7482 => x"96",     7483 => x"96",     7484 => x"95",     7485 => x"95",     7486 => x"94",     7487 => x"94", 
    7488 => x"94",     7489 => x"94",     7490 => x"94",     7491 => x"94",     7492 => x"93",     7493 => x"93",     7494 => x"92",     7495 => x"92", 
    7496 => x"91",     7497 => x"90",     7498 => x"8F",     7499 => x"90",     7500 => x"8D",     7501 => x"8C",     7502 => x"8B",     7503 => x"8B", 
    7504 => x"8C",     7505 => x"87",     7506 => x"87",     7507 => x"86",     7508 => x"88",     7509 => x"86",     7510 => x"85",     7511 => x"89", 
    7512 => x"89",     7513 => x"89",     7514 => x"89",     7515 => x"89",     7516 => x"89",     7517 => x"89",     7518 => x"89",     7519 => x"89", 
    7520 => x"89",     7521 => x"89",     7522 => x"89",     7523 => x"89",     7524 => x"89",     7525 => x"89",     7526 => x"89",     7527 => x"89", 
    7528 => x"89",     7529 => x"89",     7530 => x"89",     7531 => x"89",     7532 => x"89",     7533 => x"89",     7534 => x"89",     7535 => x"89", 
    7536 => x"89",     7537 => x"89",     7538 => x"89",     7539 => x"89",     7540 => x"89",     7541 => x"89",     7542 => x"89",     7543 => x"89", 
    7544 => x"89",     7545 => x"89",     7546 => x"89",     7547 => x"89",     7548 => x"89",     7549 => x"89",     7550 => x"89",     7551 => x"89", 
    7552 => x"89",     7553 => x"89",     7554 => x"89",     7555 => x"89",     7556 => x"89",     7557 => x"89",     7558 => x"89",     7559 => x"89", 
    7560 => x"89",     7561 => x"89",     7562 => x"89",     7563 => x"89",     7564 => x"89",     7565 => x"89",     7566 => x"89",     7567 => x"89", 
    7568 => x"89",     7569 => x"89",     7570 => x"89",     7571 => x"89",     7572 => x"89",     7573 => x"89",     7574 => x"89",     7575 => x"89", 
    7576 => x"89",     7577 => x"89",     7578 => x"89",     7579 => x"89",     7580 => x"89",     7581 => x"89",     7582 => x"89",     7583 => x"89", 
    7584 => x"89",     7585 => x"89",     7586 => x"89",     7587 => x"89",     7588 => x"89",     7589 => x"89",     7590 => x"89",     7591 => x"89", 
    7592 => x"89",     7593 => x"89",     7594 => x"89",     7595 => x"89",     7596 => x"89",     7597 => x"89",     7598 => x"89",     7599 => x"89", 
    7600 => x"89",     7601 => x"89",     7602 => x"89",     7603 => x"89",     7604 => x"89",     7605 => x"89",     7606 => x"89",     7607 => x"89", 
    7608 => x"89",     7609 => x"89",     7610 => x"89",     7611 => x"89",     7612 => x"89",     7613 => x"89",     7614 => x"89",     7615 => x"89", 
    7616 => x"89",     7617 => x"89",     7618 => x"89",     7619 => x"89",     7620 => x"89",     7621 => x"89",     7622 => x"89",     7623 => x"89", 
    7624 => x"89",     7625 => x"89",     7626 => x"89",     7627 => x"89",     7628 => x"89",     7629 => x"89",     7630 => x"89",     7631 => x"89", 
    7632 => x"89",     7633 => x"89",     7634 => x"89",     7635 => x"89",     7636 => x"89"
);


    signal sLUT : sine_table_t := (
    0 => x"80", 1 => x"86", 2 => x"8c", 3 => x"92", 4 => x"98", 5 => x"9e", 6 => x"a5", 7 => x"aa",
    8 => x"b0", 9 => x"b6", 10 => x"bc", 11 => x"c1", 12 => x"c6", 13 => x"cb", 14 => x"d0", 15 => x"d5",
    16 => x"da", 17 => x"de", 18 => x"e2", 19 => x"e6", 20 => x"ea", 21 => x"ed", 22 => x"f0", 23 => x"f3",
    24 => x"f5", 25 => x"f8", 26 => x"fa", 27 => x"fb", 28 => x"fd", 29 => x"fe", 30 => x"fe", 31 => x"ff",
    32 => x"ff", 33 => x"ff", 34 => x"fe", 35 => x"fe", 36 => x"fd", 37 => x"fb", 38 => x"fa", 39 => x"f8",
    40 => x"f5", 41 => x"f3", 42 => x"f0", 43 => x"ed", 44 => x"ea", 45 => x"e6", 46 => x"e2", 47 => x"de",
    48 => x"da", 49 => x"d5", 50 => x"d0", 51 => x"cb", 52 => x"c6", 53 => x"c1", 54 => x"bc", 55 => x"b6",
    56 => x"b0", 57 => x"aa", 58 => x"a5", 59 => x"9e", 60 => x"98", 61 => x"92", 62 => x"8c", 63 => x"86",
    64 => x"80", 65 => x"79", 66 => x"73", 67 => x"6d", 68 => x"67", 69 => x"61", 70 => x"5a", 71 => x"55",
    72 => x"4f", 73 => x"49", 74 => x"43", 75 => x"3e", 76 => x"39", 77 => x"34", 78 => x"2f", 79 => x"2a",
    80 => x"25", 81 => x"21", 82 => x"1d", 83 => x"19", 84 => x"15", 85 => x"12", 86 => x"0f", 87 => x"0c",
    88 => x"0a", 89 => x"07", 90 => x"05", 91 => x"04", 92 => x"02", 93 => x"01", 94 => x"01", 95 => x"00",
    96 => x"00", 97 => x"00", 98 => x"01", 99 => x"01", 100 => x"02", 101 => x"04", 102 => x"05", 103 => x"07",
    104 => x"0a", 105 => x"0c", 106 => x"0f", 107 => x"12", 108 => x"15", 109 => x"19", 110 => x"1d", 111 => x"21",
    112 => x"25", 113 => x"2a", 114 => x"2f", 115 => x"34", 116 => x"39", 117 => x"3e", 118 => x"43", 119 => x"49",
    120 => x"4f", 121 => x"55", 122 => x"5a", 123 => x"61", 124 => x"67", 125 => x"6d", 126 => x"73", 127 => x"79"
    );


    signal vwoopLUT : vwoop_table_t := (
    0 => x"50",     1 => x"50",     2 => x"50",     3 => x"50",     4 => x"50",     5 => x"50",     6 => x"50",     7 => x"50", 
    8 => x"50",     9 => x"50",     10 => x"50",     11 => x"50",     12 => x"50",     13 => x"50",     14 => x"50",     15 => x"50", 
    16 => x"50",     17 => x"50",     18 => x"50",     19 => x"50",     20 => x"50",     21 => x"50",     22 => x"50",     23 => x"50", 
    24 => x"50",     25 => x"50",     26 => x"50",     27 => x"50",     28 => x"50",     29 => x"50",     30 => x"50",     31 => x"50", 
    32 => x"50",     33 => x"50",     34 => x"50",     35 => x"50",     36 => x"50",     37 => x"50",     38 => x"50",     39 => x"50", 
    40 => x"50",     41 => x"50",     42 => x"50",     43 => x"50",     44 => x"50",     45 => x"50",     46 => x"50",     47 => x"50", 
    48 => x"50",     49 => x"50",     50 => x"50",     51 => x"50",     52 => x"50",     53 => x"50",     54 => x"50",     55 => x"50", 
    56 => x"50",     57 => x"00",     58 => x"00",     59 => x"00",     60 => x"00",     61 => x"00",     62 => x"00",     63 => x"00", 
    64 => x"00",     65 => x"00",     66 => x"00",     67 => x"00",     68 => x"00",     69 => x"00",     70 => x"00",     71 => x"00", 
    72 => x"00",     73 => x"00",     74 => x"00",     75 => x"00",     76 => x"00",     77 => x"00",     78 => x"00",     79 => x"00", 
    80 => x"00",     81 => x"00",     82 => x"00",     83 => x"00",     84 => x"00",     85 => x"00",     86 => x"00",     87 => x"00", 
    88 => x"00",     89 => x"00",     90 => x"00",     91 => x"00",     92 => x"00",     93 => x"00",     94 => x"00",     95 => x"00", 
    96 => x"00",     97 => x"00",     98 => x"00",     99 => x"00",     100 => x"00",     101 => x"00",     102 => x"50",     103 => x"50", 
    104 => x"50",     105 => x"50",     106 => x"50",     107 => x"50",     108 => x"50",     109 => x"50",     110 => x"50",     111 => x"50", 
    112 => x"50",     113 => x"50",     114 => x"50",     115 => x"50",     116 => x"50",     117 => x"50",     118 => x"50",     119 => x"50", 
    120 => x"50",     121 => x"50",     122 => x"50",     123 => x"50",     124 => x"50",     125 => x"50",     126 => x"50",     127 => x"50", 
    128 => x"50",     129 => x"50",     130 => x"50",     131 => x"50",     132 => x"50",     133 => x"50",     134 => x"50",     135 => x"50", 
    136 => x"50",     137 => x"50",     138 => x"50",     139 => x"50",     140 => x"00",     141 => x"00",     142 => x"00",     143 => x"00", 
    144 => x"00",     145 => x"00",     146 => x"00",     147 => x"00",     148 => x"00",     149 => x"00",     150 => x"00",     151 => x"00", 
    152 => x"00",     153 => x"00",     154 => x"00",     155 => x"00",     156 => x"00",     157 => x"00",     158 => x"00",     159 => x"00", 
    160 => x"00",     161 => x"00",     162 => x"00",     163 => x"00",     164 => x"00",     165 => x"00",     166 => x"00",     167 => x"00", 
    168 => x"00",     169 => x"00",     170 => x"00",     171 => x"00",     172 => x"00",     173 => x"00",     174 => x"50",     175 => x"50", 
    176 => x"50",     177 => x"50",     178 => x"50",     179 => x"50",     180 => x"50",     181 => x"50",     182 => x"50",     183 => x"50", 
    184 => x"50",     185 => x"50",     186 => x"50",     187 => x"50",     188 => x"50",     189 => x"50",     190 => x"50",     191 => x"50", 
    192 => x"50",     193 => x"50",     194 => x"50",     195 => x"50",     196 => x"50",     197 => x"50",     198 => x"50",     199 => x"50", 
    200 => x"50",     201 => x"50",     202 => x"50",     203 => x"50",     204 => x"50",     205 => x"00",     206 => x"00",     207 => x"00", 
    208 => x"00",     209 => x"00",     210 => x"00",     211 => x"00",     212 => x"00",     213 => x"00",     214 => x"00",     215 => x"00", 
    216 => x"00",     217 => x"00",     218 => x"00",     219 => x"00",     220 => x"00",     221 => x"00",     222 => x"00",     223 => x"00", 
    224 => x"00",     225 => x"00",     226 => x"00",     227 => x"00",     228 => x"00",     229 => x"00",     230 => x"00",     231 => x"00", 
    232 => x"00",     233 => x"50",     234 => x"50",     235 => x"50",     236 => x"50",     237 => x"50",     238 => x"50",     239 => x"50", 
    240 => x"50",     241 => x"50",     242 => x"50",     243 => x"50",     244 => x"50",     245 => x"50",     246 => x"50",     247 => x"50", 
    248 => x"50",     249 => x"50",     250 => x"50",     251 => x"50",     252 => x"50",     253 => x"50",     254 => x"50",     255 => x"50", 
    256 => x"50",     257 => x"50",     258 => x"50",     259 => x"50",     260 => x"00",     261 => x"00",     262 => x"00",     263 => x"00", 
    264 => x"00",     265 => x"00",     266 => x"00",     267 => x"00",     268 => x"00",     269 => x"00",     270 => x"00",     271 => x"00", 
    272 => x"00",     273 => x"00",     274 => x"00",     275 => x"00",     276 => x"00",     277 => x"00",     278 => x"00",     279 => x"00", 
    280 => x"00",     281 => x"00",     282 => x"00",     283 => x"00",     284 => x"00",     285 => x"50",     286 => x"50",     287 => x"50", 
    288 => x"50",     289 => x"50",     290 => x"50",     291 => x"50",     292 => x"50",     293 => x"50",     294 => x"50",     295 => x"50", 
    296 => x"50",     297 => x"50",     298 => x"50",     299 => x"50",     300 => x"50",     301 => x"50",     302 => x"50",     303 => x"50", 
    304 => x"50",     305 => x"50",     306 => x"50",     307 => x"50",     308 => x"00",     309 => x"00",     310 => x"00",     311 => x"00", 
    312 => x"00",     313 => x"00",     314 => x"00",     315 => x"00",     316 => x"00",     317 => x"00",     318 => x"00",     319 => x"00", 
    320 => x"00",     321 => x"00",     322 => x"00",     323 => x"00",     324 => x"00",     325 => x"00",     326 => x"00",     327 => x"00", 
    328 => x"00",     329 => x"00",     330 => x"00",     331 => x"50",     332 => x"50",     333 => x"50",     334 => x"50",     335 => x"50", 
    336 => x"50",     337 => x"50",     338 => x"50",     339 => x"50",     340 => x"50",     341 => x"50",     342 => x"50",     343 => x"50", 
    344 => x"50",     345 => x"50",     346 => x"50",     347 => x"50",     348 => x"50",     349 => x"50",     350 => x"50",     351 => x"50", 
    352 => x"00",     353 => x"00",     354 => x"00",     355 => x"00",     356 => x"00",     357 => x"00",     358 => x"00",     359 => x"00", 
    360 => x"00",     361 => x"00",     362 => x"00",     363 => x"00",     364 => x"00",     365 => x"00",     366 => x"00",     367 => x"00", 
    368 => x"00",     369 => x"00",     370 => x"00",     371 => x"00",     372 => x"00",     373 => x"50",     374 => x"50",     375 => x"50", 
    376 => x"50",     377 => x"50",     378 => x"50",     379 => x"50",     380 => x"50",     381 => x"50",     382 => x"50",     383 => x"50", 
    384 => x"50",     385 => x"50",     386 => x"50",     387 => x"50",     388 => x"50",     389 => x"50",     390 => x"50",     391 => x"50", 
    392 => x"50",     393 => x"00",     394 => x"00",     395 => x"00",     396 => x"00",     397 => x"00",     398 => x"00",     399 => x"00", 
    400 => x"00",     401 => x"00",     402 => x"00",     403 => x"00",     404 => x"00",     405 => x"00",     406 => x"00",     407 => x"00", 
    408 => x"00",     409 => x"00",     410 => x"00",     411 => x"00",     412 => x"50",     413 => x"50",     414 => x"50",     415 => x"50", 
    416 => x"50",     417 => x"50",     418 => x"50",     419 => x"50",     420 => x"50",     421 => x"50",     422 => x"50",     423 => x"50", 
    424 => x"50",     425 => x"50",     426 => x"50",     427 => x"50",     428 => x"50",     429 => x"50",     430 => x"00",     431 => x"00", 
    432 => x"00",     433 => x"00",     434 => x"00",     435 => x"00",     436 => x"00",     437 => x"00",     438 => x"00",     439 => x"00", 
    440 => x"00",     441 => x"00",     442 => x"00",     443 => x"00",     444 => x"00",     445 => x"00",     446 => x"00",     447 => x"00", 
    448 => x"50",     449 => x"50",     450 => x"50",     451 => x"50",     452 => x"50",     453 => x"50",     454 => x"50",     455 => x"50", 
    456 => x"50",     457 => x"50",     458 => x"50",     459 => x"50",     460 => x"50",     461 => x"50",     462 => x"50",     463 => x"50", 
    464 => x"50",     465 => x"50",     466 => x"00",     467 => x"00",     468 => x"00",     469 => x"00",     470 => x"00",     471 => x"00", 
    472 => x"00",     473 => x"00",     474 => x"00",     475 => x"00",     476 => x"00",     477 => x"00",     478 => x"00",     479 => x"00", 
    480 => x"00",     481 => x"00",     482 => x"00",     483 => x"50",     484 => x"50",     485 => x"50",     486 => x"50",     487 => x"50", 
    488 => x"50",     489 => x"50",     490 => x"50",     491 => x"50",     492 => x"50",     493 => x"50",     494 => x"50",     495 => x"50", 
    496 => x"50",     497 => x"50",     498 => x"50",     499 => x"00",     500 => x"00",     501 => x"00",     502 => x"00",     503 => x"00", 
    504 => x"00",     505 => x"00",     506 => x"00",     507 => x"00",     508 => x"00",     509 => x"00",     510 => x"00",     511 => x"00", 
    512 => x"00",     513 => x"00",     514 => x"00",     515 => x"00",     516 => x"50",     517 => x"50",     518 => x"50",     519 => x"50", 
    520 => x"50",     521 => x"50",     522 => x"50",     523 => x"50",     524 => x"50",     525 => x"50",     526 => x"50",     527 => x"50", 
    528 => x"50",     529 => x"50",     530 => x"50",     531 => x"00",     532 => x"00",     533 => x"00",     534 => x"00",     535 => x"00", 
    536 => x"00",     537 => x"00",     538 => x"00",     539 => x"00",     540 => x"00",     541 => x"00",     542 => x"00",     543 => x"00", 
    544 => x"00",     545 => x"00",     546 => x"00",     547 => x"50",     548 => x"50",     549 => x"50",     550 => x"50",     551 => x"50", 
    552 => x"50",     553 => x"50",     554 => x"50",     555 => x"50",     556 => x"50",     557 => x"50",     558 => x"50",     559 => x"50", 
    560 => x"50",     561 => x"50",     562 => x"00",     563 => x"00",     564 => x"00",     565 => x"00",     566 => x"00",     567 => x"00", 
    568 => x"00",     569 => x"00",     570 => x"00",     571 => x"00",     572 => x"00",     573 => x"00",     574 => x"00",     575 => x"00", 
    576 => x"00",     577 => x"50",     578 => x"50",     579 => x"50",     580 => x"50",     581 => x"50",     582 => x"50",     583 => x"50", 
    584 => x"50",     585 => x"50",     586 => x"50",     587 => x"50",     588 => x"50",     589 => x"50",     590 => x"50",     591 => x"00", 
    592 => x"00",     593 => x"00",     594 => x"00",     595 => x"00",     596 => x"00",     597 => x"00",     598 => x"00",     599 => x"00", 
    600 => x"00",     601 => x"00",     602 => x"00",     603 => x"00",     604 => x"00",     605 => x"50",     606 => x"50",     607 => x"50", 
    608 => x"50",     609 => x"50",     610 => x"50",     611 => x"50",     612 => x"50",     613 => x"50",     614 => x"50",     615 => x"50", 
    616 => x"50",     617 => x"50",     618 => x"50",     619 => x"00",     620 => x"00",     621 => x"00",     622 => x"00",     623 => x"00", 
    624 => x"00",     625 => x"00",     626 => x"00",     627 => x"00",     628 => x"00",     629 => x"00",     630 => x"00",     631 => x"00", 
    632 => x"00",     633 => x"50",     634 => x"50",     635 => x"50",     636 => x"50",     637 => x"50",     638 => x"50",     639 => x"50", 
    640 => x"50",     641 => x"50",     642 => x"50",     643 => x"50",     644 => x"50",     645 => x"50",     646 => x"50",     647 => x"00", 
    648 => x"00",     649 => x"00",     650 => x"00",     651 => x"00",     652 => x"00",     653 => x"00",     654 => x"00",     655 => x"00", 
    656 => x"00",     657 => x"00",     658 => x"00",     659 => x"00",     660 => x"50",     661 => x"50",     662 => x"50",     663 => x"50", 
    664 => x"50",     665 => x"50",     666 => x"50",     667 => x"50",     668 => x"50",     669 => x"50",     670 => x"50",     671 => x"50", 
    672 => x"50",     673 => x"00",     674 => x"00",     675 => x"00",     676 => x"00",     677 => x"00",     678 => x"00",     679 => x"00", 
    680 => x"00",     681 => x"00",     682 => x"00",     683 => x"00",     684 => x"00",     685 => x"00",     686 => x"50",     687 => x"50", 
    688 => x"50",     689 => x"50",     690 => x"50",     691 => x"50",     692 => x"50",     693 => x"50",     694 => x"50",     695 => x"50", 
    696 => x"50",     697 => x"50",     698 => x"00",     699 => x"00",     700 => x"00",     701 => x"00",     702 => x"00",     703 => x"00", 
    704 => x"00",     705 => x"00",     706 => x"00",     707 => x"00",     708 => x"00",     709 => x"00",     710 => x"00",     711 => x"50", 
    712 => x"50",     713 => x"50",     714 => x"50",     715 => x"50",     716 => x"50",     717 => x"50",     718 => x"50",     719 => x"50", 
    720 => x"50",     721 => x"50",     722 => x"50",     723 => x"00",     724 => x"00",     725 => x"00",     726 => x"00",     727 => x"00", 
    728 => x"00",     729 => x"00",     730 => x"00",     731 => x"00",     732 => x"00",     733 => x"00",     734 => x"00",     735 => x"50", 
    736 => x"50",     737 => x"50",     738 => x"50",     739 => x"50",     740 => x"50",     741 => x"50",     742 => x"50",     743 => x"50", 
    744 => x"50",     745 => x"50",     746 => x"50",     747 => x"00",     748 => x"00",     749 => x"00",     750 => x"00",     751 => x"00", 
    752 => x"00",     753 => x"00",     754 => x"00",     755 => x"00",     756 => x"00",     757 => x"00",     758 => x"00",     759 => x"50", 
    760 => x"50",     761 => x"50",     762 => x"50",     763 => x"50",     764 => x"50",     765 => x"50",     766 => x"50",     767 => x"50", 
    768 => x"50",     769 => x"50",     770 => x"50",     771 => x"00",     772 => x"00",     773 => x"00",     774 => x"00",     775 => x"00", 
    776 => x"00",     777 => x"00",     778 => x"00",     779 => x"00",     780 => x"00",     781 => x"00",     782 => x"50",     783 => x"50", 
    784 => x"50",     785 => x"50",     786 => x"50",     787 => x"50",     788 => x"50",     789 => x"50",     790 => x"50",     791 => x"50", 
    792 => x"50",     793 => x"50",     794 => x"00",     795 => x"00",     796 => x"00",     797 => x"00",     798 => x"00",     799 => x"00", 
    800 => x"00",     801 => x"00",     802 => x"00",     803 => x"00",     804 => x"00",     805 => x"50",     806 => x"50",     807 => x"50", 
    808 => x"50",     809 => x"50",     810 => x"50",     811 => x"50",     812 => x"50",     813 => x"50",     814 => x"50",     815 => x"50", 
    816 => x"00",     817 => x"00",     818 => x"00",     819 => x"00",     820 => x"00",     821 => x"00",     822 => x"00",     823 => x"00", 
    824 => x"00",     825 => x"00",     826 => x"00",     827 => x"50",     828 => x"50",     829 => x"50",     830 => x"50",     831 => x"50", 
    832 => x"50",     833 => x"50",     834 => x"50",     835 => x"50",     836 => x"50",     837 => x"50",     838 => x"00",     839 => x"00", 
    840 => x"00",     841 => x"00",     842 => x"00",     843 => x"00",     844 => x"00",     845 => x"00",     846 => x"00",     847 => x"00", 
    848 => x"00",     849 => x"50",     850 => x"50",     851 => x"50",     852 => x"50",     853 => x"50",     854 => x"50",     855 => x"50", 
    856 => x"50",     857 => x"50",     858 => x"50",     859 => x"00",     860 => x"00",     861 => x"00",     862 => x"00",     863 => x"00", 
    864 => x"00",     865 => x"00",     866 => x"00",     867 => x"00",     868 => x"00",     869 => x"00",     870 => x"50",     871 => x"50", 
    872 => x"50",     873 => x"50",     874 => x"50",     875 => x"50",     876 => x"50",     877 => x"50",     878 => x"50",     879 => x"50", 
    880 => x"00",     881 => x"00",     882 => x"00",     883 => x"00",     884 => x"00",     885 => x"00",     886 => x"00",     887 => x"00", 
    888 => x"00",     889 => x"00",     890 => x"00",     891 => x"50",     892 => x"50",     893 => x"50",     894 => x"50",     895 => x"50", 
    896 => x"50",     897 => x"50",     898 => x"50",     899 => x"50",     900 => x"50",     901 => x"00",     902 => x"00",     903 => x"00", 
    904 => x"00",     905 => x"00",     906 => x"00",     907 => x"00",     908 => x"00",     909 => x"00",     910 => x"00",     911 => x"50", 
    912 => x"50",     913 => x"50",     914 => x"50",     915 => x"50",     916 => x"50",     917 => x"50",     918 => x"50",     919 => x"50", 
    920 => x"50",     921 => x"00",     922 => x"00",     923 => x"00",     924 => x"00",     925 => x"00",     926 => x"00",     927 => x"00", 
    928 => x"00",     929 => x"00",     930 => x"00",     931 => x"50",     932 => x"50",     933 => x"50",     934 => x"50",     935 => x"50", 
    936 => x"50",     937 => x"50",     938 => x"50",     939 => x"50",     940 => x"50",     941 => x"00",     942 => x"00",     943 => x"00", 
    944 => x"00",     945 => x"00",     946 => x"00",     947 => x"00",     948 => x"00",     949 => x"00",     950 => x"00",     951 => x"50", 
    952 => x"50",     953 => x"50",     954 => x"50",     955 => x"50",     956 => x"50",     957 => x"50",     958 => x"50",     959 => x"50", 
    960 => x"00",     961 => x"00",     962 => x"00",     963 => x"00",     964 => x"00",     965 => x"00",     966 => x"00",     967 => x"00", 
    968 => x"00",     969 => x"00",     970 => x"50",     971 => x"50",     972 => x"50",     973 => x"50",     974 => x"50",     975 => x"50", 
    976 => x"50",     977 => x"50",     978 => x"50",     979 => x"00",     980 => x"00",     981 => x"00",     982 => x"00",     983 => x"00", 
    984 => x"00",     985 => x"00",     986 => x"00",     987 => x"00",     988 => x"00",     989 => x"50",     990 => x"50",     991 => x"50", 
    992 => x"50",     993 => x"50",     994 => x"50",     995 => x"50",     996 => x"50",     997 => x"50",     998 => x"00",     999 => x"00", 
    1000 => x"00",     1001 => x"00",     1002 => x"00",     1003 => x"00",     1004 => x"00",     1005 => x"00",     1006 => x"00",     1007 => x"50", 
    1008 => x"50",     1009 => x"50",     1010 => x"50",     1011 => x"50",     1012 => x"50",     1013 => x"50",     1014 => x"50",     1015 => x"50", 
    1016 => x"50",     1017 => x"00",     1018 => x"00",     1019 => x"00",     1020 => x"00",     1021 => x"00",     1022 => x"00",     1023 => x"00", 
    1024 => x"00",     1025 => x"00",     1026 => x"50",     1027 => x"50",     1028 => x"50",     1029 => x"50",     1030 => x"50",     1031 => x"50", 
    1032 => x"50",     1033 => x"50",     1034 => x"50",     1035 => x"00",     1036 => x"00",     1037 => x"00",     1038 => x"00",     1039 => x"00", 
    1040 => x"00",     1041 => x"00",     1042 => x"00",     1043 => x"00",     1044 => x"50",     1045 => x"50",     1046 => x"50",     1047 => x"50", 
    1048 => x"50",     1049 => x"50",     1050 => x"50",     1051 => x"50",     1052 => x"50",     1053 => x"00",     1054 => x"00",     1055 => x"00", 
    1056 => x"00",     1057 => x"00",     1058 => x"00",     1059 => x"00",     1060 => x"00",     1061 => x"00",     1062 => x"50",     1063 => x"50", 
    1064 => x"50",     1065 => x"50",     1066 => x"50",     1067 => x"50",     1068 => x"50",     1069 => x"50",     1070 => x"00",     1071 => x"00", 
    1072 => x"00",     1073 => x"00",     1074 => x"00",     1075 => x"00",     1076 => x"00",     1077 => x"00",     1078 => x"00",     1079 => x"50", 
    1080 => x"50",     1081 => x"50",     1082 => x"50",     1083 => x"50",     1084 => x"50",     1085 => x"50",     1086 => x"50",     1087 => x"50", 
    1088 => x"00",     1089 => x"00",     1090 => x"00",     1091 => x"00",     1092 => x"00",     1093 => x"00",     1094 => x"00",     1095 => x"00", 
    1096 => x"00",     1097 => x"50",     1098 => x"50",     1099 => x"50",     1100 => x"50",     1101 => x"50",     1102 => x"50",     1103 => x"50", 
    1104 => x"50",     1105 => x"00",     1106 => x"00",     1107 => x"00",     1108 => x"00",     1109 => x"00",     1110 => x"00",     1111 => x"00", 
    1112 => x"00",     1113 => x"00",     1114 => x"50",     1115 => x"50",     1116 => x"50",     1117 => x"50",     1118 => x"50",     1119 => x"50", 
    1120 => x"50",     1121 => x"50",     1122 => x"00",     1123 => x"00",     1124 => x"00",     1125 => x"00",     1126 => x"00",     1127 => x"00", 
    1128 => x"00",     1129 => x"00",     1130 => x"50",     1131 => x"50",     1132 => x"50",     1133 => x"50",     1134 => x"50",     1135 => x"50", 
    1136 => x"50",     1137 => x"50",     1138 => x"50",     1139 => x"00",     1140 => x"00",     1141 => x"00",     1142 => x"00",     1143 => x"00", 
    1144 => x"00",     1145 => x"00",     1146 => x"00",     1147 => x"50",     1148 => x"50",     1149 => x"50",     1150 => x"50",     1151 => x"50", 
    1152 => x"50",     1153 => x"50",     1154 => x"50",     1155 => x"00",     1156 => x"00",     1157 => x"00",     1158 => x"00",     1159 => x"00", 
    1160 => x"00",     1161 => x"00",     1162 => x"00",     1163 => x"50",     1164 => x"50",     1165 => x"50",     1166 => x"50",     1167 => x"50", 
    1168 => x"50",     1169 => x"50",     1170 => x"50",     1171 => x"50",     1172 => x"00",     1173 => x"00",     1174 => x"00",     1175 => x"00", 
    1176 => x"00",     1177 => x"00",     1178 => x"00",     1179 => x"00",     1180 => x"50",     1181 => x"50",     1182 => x"50",     1183 => x"50", 
    1184 => x"50",     1185 => x"50",     1186 => x"50",     1187 => x"50",     1188 => x"00",     1189 => x"00",     1190 => x"00",     1191 => x"00", 
    1192 => x"00",     1193 => x"00",     1194 => x"00",     1195 => x"00",     1196 => x"50",     1197 => x"50",     1198 => x"50",     1199 => x"50", 
    1200 => x"50",     1201 => x"50",     1202 => x"50",     1203 => x"50",     1204 => x"00",     1205 => x"00",     1206 => x"00",     1207 => x"00", 
    1208 => x"00",     1209 => x"00",     1210 => x"00",     1211 => x"00",     1212 => x"50",     1213 => x"50",     1214 => x"50",     1215 => x"50", 
    1216 => x"50",     1217 => x"50",     1218 => x"50",     1219 => x"00",     1220 => x"00",     1221 => x"00",     1222 => x"00",     1223 => x"00", 
    1224 => x"00",     1225 => x"00",     1226 => x"00",     1227 => x"50",     1228 => x"50",     1229 => x"50",     1230 => x"50",     1231 => x"50", 
    1232 => x"50",     1233 => x"50",     1234 => x"50",     1235 => x"00",     1236 => x"00",     1237 => x"00",     1238 => x"00",     1239 => x"00", 
    1240 => x"00",     1241 => x"00",     1242 => x"00",     1243 => x"50",     1244 => x"50",     1245 => x"50",     1246 => x"50",     1247 => x"50", 
    1248 => x"50",     1249 => x"50",     1250 => x"00",     1251 => x"00",     1252 => x"00",     1253 => x"00",     1254 => x"00",     1255 => x"00", 
    1256 => x"00",     1257 => x"00",     1258 => x"50",     1259 => x"50",     1260 => x"50",     1261 => x"50",     1262 => x"50",     1263 => x"50", 
    1264 => x"50",     1265 => x"50",     1266 => x"00",     1267 => x"00",     1268 => x"00",     1269 => x"00",     1270 => x"00",     1271 => x"00", 
    1272 => x"00",     1273 => x"50",     1274 => x"50",     1275 => x"50",     1276 => x"50",     1277 => x"50",     1278 => x"50",     1279 => x"50", 
    1280 => x"50",     1281 => x"00",     1282 => x"00",     1283 => x"00",     1284 => x"00",     1285 => x"00",     1286 => x"00",     1287 => x"00", 
    1288 => x"50",     1289 => x"50",     1290 => x"50",     1291 => x"50",     1292 => x"50",     1293 => x"50",     1294 => x"50",     1295 => x"50", 
    1296 => x"00",     1297 => x"00",     1298 => x"00",     1299 => x"00",     1300 => x"00",     1301 => x"00",     1302 => x"00",     1303 => x"50", 
    1304 => x"50",     1305 => x"50",     1306 => x"50",     1307 => x"50",     1308 => x"50",     1309 => x"50",     1310 => x"00",     1311 => x"00", 
    1312 => x"00",     1313 => x"00",     1314 => x"00",     1315 => x"00",     1316 => x"00",     1317 => x"00",     1318 => x"50",     1319 => x"50", 
    1320 => x"50",     1321 => x"50",     1322 => x"50",     1323 => x"50",     1324 => x"50",     1325 => x"00",     1326 => x"00",     1327 => x"00", 
    1328 => x"00",     1329 => x"00",     1330 => x"00",     1331 => x"00",     1332 => x"50",     1333 => x"50",     1334 => x"50",     1335 => x"50", 
    1336 => x"50",     1337 => x"50",     1338 => x"50",     1339 => x"00",     1340 => x"00",     1341 => x"00",     1342 => x"00",     1343 => x"00", 
    1344 => x"00",     1345 => x"00",     1346 => x"00",     1347 => x"50",     1348 => x"50",     1349 => x"50",     1350 => x"50",     1351 => x"50", 
    1352 => x"50",     1353 => x"50",     1354 => x"00",     1355 => x"00",     1356 => x"00",     1357 => x"00",     1358 => x"00",     1359 => x"00", 
    1360 => x"00",     1361 => x"50",     1362 => x"50",     1363 => x"50",     1364 => x"50",     1365 => x"50",     1366 => x"50",     1367 => x"50", 
    1368 => x"00",     1369 => x"00",     1370 => x"00",     1371 => x"00",     1372 => x"00",     1373 => x"00",     1374 => x"00",     1375 => x"50", 
    1376 => x"50",     1377 => x"50",     1378 => x"50",     1379 => x"50",     1380 => x"50",     1381 => x"50",     1382 => x"00",     1383 => x"00", 
    1384 => x"00",     1385 => x"00",     1386 => x"00",     1387 => x"00",     1388 => x"00",     1389 => x"50",     1390 => x"50",     1391 => x"50", 
    1392 => x"50",     1393 => x"50",     1394 => x"50",     1395 => x"50",     1396 => x"00",     1397 => x"00",     1398 => x"00",     1399 => x"00", 
    1400 => x"00",     1401 => x"00",     1402 => x"00",     1403 => x"50",     1404 => x"50",     1405 => x"50",     1406 => x"50",     1407 => x"50", 
    1408 => x"50",     1409 => x"50",     1410 => x"00",     1411 => x"00",     1412 => x"00",     1413 => x"00",     1414 => x"00",     1415 => x"00", 
    1416 => x"00",     1417 => x"50",     1418 => x"50",     1419 => x"50",     1420 => x"50",     1421 => x"50",     1422 => x"50",     1423 => x"50", 
    1424 => x"00",     1425 => x"00",     1426 => x"00",     1427 => x"00",     1428 => x"00",     1429 => x"00",     1430 => x"50",     1431 => x"50", 
    1432 => x"50",     1433 => x"50",     1434 => x"50",     1435 => x"50",     1436 => x"50",     1437 => x"00",     1438 => x"00",     1439 => x"00", 
    1440 => x"00",     1441 => x"00",     1442 => x"00",     1443 => x"00",     1444 => x"50",     1445 => x"50",     1446 => x"50",     1447 => x"50", 
    1448 => x"50",     1449 => x"50",     1450 => x"50",     1451 => x"00",     1452 => x"00",     1453 => x"00",     1454 => x"00",     1455 => x"00", 
    1456 => x"00",     1457 => x"50",     1458 => x"50",     1459 => x"50",     1460 => x"50",     1461 => x"50",     1462 => x"50",     1463 => x"50", 
    1464 => x"00",     1465 => x"00",     1466 => x"00",     1467 => x"00",     1468 => x"00",     1469 => x"00",     1470 => x"00",     1471 => x"50", 
    1472 => x"50",     1473 => x"50",     1474 => x"50",     1475 => x"50",     1476 => x"50",     1477 => x"00",     1478 => x"00",     1479 => x"00", 
    1480 => x"00",     1481 => x"00",     1482 => x"00",     1483 => x"00",     1484 => x"50",     1485 => x"50",     1486 => x"50",     1487 => x"50", 
    1488 => x"50",     1489 => x"50",     1490 => x"00",     1491 => x"00",     1492 => x"00",     1493 => x"00",     1494 => x"00",     1495 => x"00", 
    1496 => x"00",     1497 => x"50",     1498 => x"50",     1499 => x"50",     1500 => x"50",     1501 => x"50",     1502 => x"50",     1503 => x"00", 
    1504 => x"00",     1505 => x"00",     1506 => x"00",     1507 => x"00",     1508 => x"00",     1509 => x"00",     1510 => x"50",     1511 => x"50", 
    1512 => x"50",     1513 => x"50",     1514 => x"50",     1515 => x"50",     1516 => x"00",     1517 => x"00",     1518 => x"00",     1519 => x"00", 
    1520 => x"00",     1521 => x"00",     1522 => x"00",     1523 => x"50",     1524 => x"50",     1525 => x"50",     1526 => x"50",     1527 => x"50", 
    1528 => x"50",     1529 => x"00",     1530 => x"00",     1531 => x"00",     1532 => x"00",     1533 => x"00",     1534 => x"00",     1535 => x"50", 
    1536 => x"50",     1537 => x"50",     1538 => x"50",     1539 => x"50",     1540 => x"50",     1541 => x"50",     1542 => x"00",     1543 => x"00", 
    1544 => x"00",     1545 => x"00",     1546 => x"00",     1547 => x"00",     1548 => x"50",     1549 => x"50",     1550 => x"50",     1551 => x"50", 
    1552 => x"50",     1553 => x"50",     1554 => x"50",     1555 => x"00",     1556 => x"00",     1557 => x"00",     1558 => x"00",     1559 => x"00", 
    1560 => x"00",     1561 => x"50",     1562 => x"50",     1563 => x"50",     1564 => x"50",     1565 => x"50",     1566 => x"50",     1567 => x"00", 
    1568 => x"00",     1569 => x"00",     1570 => x"00",     1571 => x"00",     1572 => x"00",     1573 => x"50",     1574 => x"50",     1575 => x"50", 
    1576 => x"50",     1577 => x"50",     1578 => x"50",     1579 => x"50",     1580 => x"00",     1581 => x"00",     1582 => x"00",     1583 => x"00", 
    1584 => x"00",     1585 => x"00",     1586 => x"50",     1587 => x"50",     1588 => x"50",     1589 => x"50",     1590 => x"50",     1591 => x"50", 
    1592 => x"00",     1593 => x"00",     1594 => x"00",     1595 => x"00",     1596 => x"00",     1597 => x"00",     1598 => x"50",     1599 => x"50", 
    1600 => x"50",     1601 => x"50",     1602 => x"50",     1603 => x"50",     1604 => x"00",     1605 => x"00",     1606 => x"00",     1607 => x"00", 
    1608 => x"00",     1609 => x"00",     1610 => x"50",     1611 => x"50",     1612 => x"50",     1613 => x"50",     1614 => x"50",     1615 => x"50", 
    1616 => x"00",     1617 => x"00",     1618 => x"00",     1619 => x"00",     1620 => x"00",     1621 => x"00",     1622 => x"50",     1623 => x"50", 
    1624 => x"50",     1625 => x"50",     1626 => x"50",     1627 => x"50",     1628 => x"00",     1629 => x"00",     1630 => x"00",     1631 => x"00", 
    1632 => x"00",     1633 => x"00",     1634 => x"00",     1635 => x"50",     1636 => x"50",     1637 => x"50",     1638 => x"50",     1639 => x"50", 
    1640 => x"50",     1641 => x"00",     1642 => x"00",     1643 => x"00",     1644 => x"00",     1645 => x"00",     1646 => x"00",     1647 => x"50", 
    1648 => x"50",     1649 => x"50",     1650 => x"50",     1651 => x"50",     1652 => x"00",     1653 => x"00",     1654 => x"00",     1655 => x"00", 
    1656 => x"00",     1657 => x"00",     1658 => x"50",     1659 => x"50",     1660 => x"50",     1661 => x"50",     1662 => x"50",     1663 => x"50", 
    1664 => x"00",     1665 => x"00",     1666 => x"00",     1667 => x"00",     1668 => x"00",     1669 => x"00",     1670 => x"50",     1671 => x"50", 
    1672 => x"50",     1673 => x"50",     1674 => x"50",     1675 => x"50",     1676 => x"00",     1677 => x"00",     1678 => x"00",     1679 => x"00", 
    1680 => x"00",     1681 => x"00",     1682 => x"50",     1683 => x"50",     1684 => x"50",     1685 => x"50",     1686 => x"50",     1687 => x"50", 
    1688 => x"00",     1689 => x"00",     1690 => x"00",     1691 => x"00",     1692 => x"00",     1693 => x"00",     1694 => x"50",     1695 => x"50", 
    1696 => x"50",     1697 => x"50",     1698 => x"50",     1699 => x"50",     1700 => x"00",     1701 => x"00",     1702 => x"00",     1703 => x"00", 
    1704 => x"00",     1705 => x"50",     1706 => x"50",     1707 => x"50",     1708 => x"50",     1709 => x"50",     1710 => x"50",     1711 => x"00", 
    1712 => x"00",     1713 => x"00",     1714 => x"00",     1715 => x"00",     1716 => x"00",     1717 => x"50",     1718 => x"50",     1719 => x"50", 
    1720 => x"50",     1721 => x"50",     1722 => x"50",     1723 => x"00",     1724 => x"00",     1725 => x"00",     1726 => x"00",     1727 => x"00", 
    1728 => x"50",     1729 => x"50",     1730 => x"50",     1731 => x"50",     1732 => x"50",     1733 => x"50",     1734 => x"00",     1735 => x"00", 
    1736 => x"00",     1737 => x"00",     1738 => x"00",     1739 => x"00",     1740 => x"50",     1741 => x"50",     1742 => x"50",     1743 => x"50", 
    1744 => x"50",     1745 => x"00",     1746 => x"00",     1747 => x"00",     1748 => x"00",     1749 => x"00",     1750 => x"00",     1751 => x"50", 
    1752 => x"50",     1753 => x"50",     1754 => x"50",     1755 => x"50",     1756 => x"50",     1757 => x"00",     1758 => x"00",     1759 => x"00", 
    1760 => x"00",     1761 => x"00",     1762 => x"50",     1763 => x"50",     1764 => x"50",     1765 => x"50",     1766 => x"50",     1767 => x"50", 
    1768 => x"00",     1769 => x"00",     1770 => x"00",     1771 => x"00",     1772 => x"00",     1773 => x"00",     1774 => x"50",     1775 => x"50", 
    1776 => x"50",     1777 => x"50",     1778 => x"50",     1779 => x"00",     1780 => x"00",     1781 => x"00",     1782 => x"00",     1783 => x"00", 
    1784 => x"00",     1785 => x"50",     1786 => x"50",     1787 => x"50",     1788 => x"50",     1789 => x"50",     1790 => x"00",     1791 => x"00", 
    1792 => x"00",     1793 => x"00",     1794 => x"00",     1795 => x"00",     1796 => x"50",     1797 => x"50",     1798 => x"50",     1799 => x"50", 
    1800 => x"50",     1801 => x"00",     1802 => x"00",     1803 => x"00",     1804 => x"00",     1805 => x"00",     1806 => x"00",     1807 => x"50", 
    1808 => x"50",     1809 => x"50",     1810 => x"50",     1811 => x"50",     1812 => x"00",     1813 => x"00",     1814 => x"00",     1815 => x"00", 
    1816 => x"00",     1817 => x"00",     1818 => x"50",     1819 => x"50",     1820 => x"50",     1821 => x"50",     1822 => x"50",     1823 => x"00", 
    1824 => x"00",     1825 => x"00",     1826 => x"00",     1827 => x"00",     1828 => x"00",     1829 => x"50",     1830 => x"50",     1831 => x"50", 
    1832 => x"50",     1833 => x"50",     1834 => x"00",     1835 => x"00",     1836 => x"00",     1837 => x"00",     1838 => x"00",     1839 => x"00", 
    1840 => x"50",     1841 => x"50",     1842 => x"50",     1843 => x"50",     1844 => x"50",     1845 => x"00",     1846 => x"00",     1847 => x"00", 
    1848 => x"00",     1849 => x"00",     1850 => x"50",     1851 => x"50",     1852 => x"50",     1853 => x"50",     1854 => x"50",     1855 => x"50", 
    1856 => x"00",     1857 => x"00",     1858 => x"00",     1859 => x"00",     1860 => x"00",     1861 => x"50",     1862 => x"50",     1863 => x"50", 
    1864 => x"50",     1865 => x"50",     1866 => x"00",     1867 => x"00",     1868 => x"00",     1869 => x"00",     1870 => x"00",     1871 => x"00", 
    1872 => x"50",     1873 => x"50",     1874 => x"50",     1875 => x"50",     1876 => x"50",     1877 => x"00",     1878 => x"00",     1879 => x"00", 
    1880 => x"00",     1881 => x"00",     1882 => x"50",     1883 => x"50",     1884 => x"50",     1885 => x"50",     1886 => x"50",     1887 => x"50", 
    1888 => x"00",     1889 => x"00",     1890 => x"00",     1891 => x"00",     1892 => x"00",     1893 => x"50",     1894 => x"50",     1895 => x"50", 
    1896 => x"50",     1897 => x"50",     1898 => x"00",     1899 => x"00",     1900 => x"00",     1901 => x"00",     1902 => x"00",     1903 => x"50", 
    1904 => x"50",     1905 => x"50",     1906 => x"50",     1907 => x"50",     1908 => x"50",     1909 => x"00",     1910 => x"00",     1911 => x"00", 
    1912 => x"00",     1913 => x"00",     1914 => x"50",     1915 => x"50",     1916 => x"50",     1917 => x"50",     1918 => x"50",     1919 => x"00", 
    1920 => x"00",     1921 => x"00",     1922 => x"00",     1923 => x"00",     1924 => x"50",     1925 => x"50",     1926 => x"50",     1927 => x"50", 
    1928 => x"50",     1929 => x"00",     1930 => x"00",     1931 => x"00",     1932 => x"00",     1933 => x"00",     1934 => x"50",     1935 => x"50", 
    1936 => x"50",     1937 => x"50",     1938 => x"50",     1939 => x"50",     1940 => x"00",     1941 => x"00",     1942 => x"00",     1943 => x"00", 
    1944 => x"00",     1945 => x"50",     1946 => x"50",     1947 => x"50",     1948 => x"50",     1949 => x"50",     1950 => x"00",     1951 => x"00", 
    1952 => x"00",     1953 => x"00",     1954 => x"00",     1955 => x"50",     1956 => x"50",     1957 => x"50",     1958 => x"50",     1959 => x"50", 
    1960 => x"00",     1961 => x"00",     1962 => x"00",     1963 => x"00",     1964 => x"00",     1965 => x"50",     1966 => x"50",     1967 => x"50", 
    1968 => x"50",     1969 => x"50",     1970 => x"00",     1971 => x"00",     1972 => x"00",     1973 => x"00",     1974 => x"00",     1975 => x"50", 
    1976 => x"50",     1977 => x"50",     1978 => x"50",     1979 => x"50",     1980 => x"00",     1981 => x"00",     1982 => x"00",     1983 => x"00", 
    1984 => x"00",     1985 => x"50",     1986 => x"50",     1987 => x"50",     1988 => x"50",     1989 => x"50",     1990 => x"00",     1991 => x"00", 
    1992 => x"00",     1993 => x"00",     1994 => x"00",     1995 => x"50",     1996 => x"50",     1997 => x"50",     1998 => x"50",     1999 => x"50"
);

signal wompLUT : womp_table_t := (
    0 => x"75",     1 => x"75",     2 => x"75",     3 => x"76",     4 => x"77",     5 => x"77",     6 => x"77",     7 => x"78", 
    8 => x"78",     9 => x"78",     10 => x"77",     11 => x"77",     12 => x"76",     13 => x"76",     14 => x"76",     15 => x"76", 
    16 => x"76",     17 => x"76",     18 => x"75",     19 => x"75",     20 => x"75",     21 => x"74",     22 => x"74",     23 => x"75", 
    24 => x"75",     25 => x"76",     26 => x"76",     27 => x"76",     28 => x"76",     29 => x"76",     30 => x"76",     31 => x"75", 
    32 => x"75",     33 => x"75",     34 => x"75",     35 => x"75",     36 => x"76",     37 => x"76",     38 => x"76",     39 => x"76", 
    40 => x"76",     41 => x"76",     42 => x"76",     43 => x"76",     44 => x"76",     45 => x"77",     46 => x"77",     47 => x"77", 
    48 => x"78",     49 => x"78",     50 => x"78",     51 => x"78",     52 => x"77",     53 => x"77",     54 => x"77",     55 => x"76", 
    56 => x"76",     57 => x"76",     58 => x"76",     59 => x"76",     60 => x"76",     61 => x"77",     62 => x"77",     63 => x"77", 
    64 => x"77",     65 => x"77",     66 => x"78",     67 => x"78",     68 => x"78",     69 => x"78",     70 => x"78",     71 => x"78", 
    72 => x"78",     73 => x"78",     74 => x"77",     75 => x"77",     76 => x"77",     77 => x"76",     78 => x"75",     79 => x"74", 
    80 => x"74",     81 => x"74",     82 => x"74",     83 => x"74",     84 => x"74",     85 => x"74",     86 => x"73",     87 => x"73", 
    88 => x"73",     89 => x"73",     90 => x"74",     91 => x"75",     92 => x"75",     93 => x"76",     94 => x"77",     95 => x"78", 
    96 => x"78",     97 => x"79",     98 => x"79",     99 => x"79",     100 => x"79",     101 => x"78",     102 => x"78",     103 => x"78", 
    104 => x"78",     105 => x"77",     106 => x"77",     107 => x"77",     108 => x"76",     109 => x"76",     110 => x"76",     111 => x"75", 
    112 => x"75",     113 => x"75",     114 => x"74",     115 => x"73",     116 => x"73",     117 => x"72",     118 => x"72",     119 => x"72", 
    120 => x"73",     121 => x"74",     122 => x"75",     123 => x"75",     124 => x"76",     125 => x"77",     126 => x"78",     127 => x"79", 
    128 => x"7A",     129 => x"7B",     130 => x"7B",     131 => x"7C",     132 => x"7C",     133 => x"7C",     134 => x"7C",     135 => x"7A", 
    136 => x"78",     137 => x"76",     138 => x"74",     139 => x"73",     140 => x"72",     141 => x"71",     142 => x"70",     143 => x"71", 
    144 => x"71",     145 => x"71",     146 => x"70",     147 => x"6F",     148 => x"71",     149 => x"73",     150 => x"75",     151 => x"75", 
    152 => x"73",     153 => x"70",     154 => x"6E",     155 => x"70",     156 => x"74",     157 => x"7A",     158 => x"81",     159 => x"86", 
    160 => x"8A",     161 => x"8B",     162 => x"8B",     163 => x"8A",     164 => x"87",     165 => x"83",     166 => x"7D",     167 => x"78", 
    168 => x"71",     169 => x"6C",     170 => x"66",     171 => x"61",     172 => x"5D",     173 => x"63",     174 => x"67",     175 => x"69", 
    176 => x"69",     177 => x"66",     178 => x"5D",     179 => x"5C",     180 => x"5E",     181 => x"65",     182 => x"72",     183 => x"80", 
    184 => x"90",     185 => x"9C",     186 => x"A3",     187 => x"A5",     188 => x"9F",     189 => x"96",     190 => x"88",     191 => x"7E", 
    192 => x"74",     193 => x"6E",     194 => x"6B",     195 => x"66",     196 => x"64",     197 => x"61",     198 => x"64",     199 => x"68", 
    200 => x"6B",     201 => x"71",     202 => x"73",     203 => x"76",     204 => x"77",     205 => x"80",     206 => x"84",     207 => x"82", 
    208 => x"7C",     209 => x"6F",     210 => x"5C",     211 => x"4F",     212 => x"48",     213 => x"4B",     214 => x"58",     215 => x"6A", 
    216 => x"7F",     217 => x"92",     218 => x"A3",     219 => x"AC",     220 => x"AF",     221 => x"AA",     222 => x"A0",     223 => x"95", 
    224 => x"87",     225 => x"7B",     226 => x"72",     227 => x"6A",     228 => x"62",     229 => x"5D",     230 => x"5B",     231 => x"5B", 
    232 => x"5E",     233 => x"63",     234 => x"68",     235 => x"6C",     236 => x"6E",     237 => x"74",     238 => x"80",     239 => x"85", 
    240 => x"85",     241 => x"7F",     242 => x"6F",     243 => x"59",     244 => x"4D",     245 => x"44",     246 => x"48",     247 => x"56", 
    248 => x"69",     249 => x"82",     250 => x"97",     251 => x"A9",     252 => x"B3",     253 => x"B5",     254 => x"AF",     255 => x"A5", 
    256 => x"9C",     257 => x"8B",     258 => x"7F",     259 => x"72",     260 => x"66",     261 => x"5D",     262 => x"57",     263 => x"56", 
    264 => x"55",     265 => x"59",     266 => x"60",     267 => x"68",     268 => x"71",     269 => x"75",     270 => x"79",     271 => x"7C", 
    272 => x"84",     273 => x"87",     274 => x"82",     275 => x"79",     276 => x"67",     277 => x"53",     278 => x"48",     279 => x"42", 
    280 => x"49",     281 => x"57",     282 => x"6D",     283 => x"86",     284 => x"9B",     285 => x"AD",     286 => x"B6",     287 => x"B9", 
    288 => x"B2",     289 => x"A7",     290 => x"9C",     291 => x"8A",     292 => x"7B",     293 => x"6E",     294 => x"63",     295 => x"59", 
    296 => x"54",     297 => x"53",     298 => x"52",     299 => x"57",     300 => x"5E",     301 => x"67",     302 => x"6E",     303 => x"74", 
    304 => x"7A",     305 => x"7F",     306 => x"8A",     307 => x"8B",     308 => x"86",     309 => x"7B",     310 => x"66",     311 => x"50", 
    312 => x"43",     313 => x"3D",     314 => x"45",     315 => x"57",     316 => x"70",     317 => x"89",     318 => x"A0",     319 => x"B3", 
    320 => x"BA",     321 => x"BB",     322 => x"B1",     323 => x"A5",     324 => x"99",     325 => x"87",     326 => x"79",     327 => x"69", 
    328 => x"5E",     329 => x"53",     330 => x"4D",     331 => x"4D",     332 => x"4D",     333 => x"55",     334 => x"5E",     335 => x"69", 
    336 => x"73",     337 => x"79",     338 => x"7D",     339 => x"80",     340 => x"8B",     341 => x"8C",     342 => x"88",     343 => x"7D", 
    344 => x"69",     345 => x"51",     346 => x"43",     347 => x"3A",     348 => x"3F",     349 => x"4E",     350 => x"66",     351 => x"82", 
    352 => x"9B",     353 => x"B2",     354 => x"BD",     355 => x"C0",     356 => x"B9",     357 => x"AC",     358 => x"9F",     359 => x"8C", 
    360 => x"7C",     361 => x"6B",     362 => x"5D",     363 => x"52",     364 => x"4B",     365 => x"4C",     366 => x"4F",     367 => x"58", 
    368 => x"62",     369 => x"6E",     370 => x"79",     371 => x"7F",     372 => x"84",     373 => x"84",     374 => x"8C",     375 => x"8F", 
    376 => x"8B",     377 => x"80",     378 => x"6E",     379 => x"53",     380 => x"3F",     381 => x"34",     382 => x"33",     383 => x"42", 
    384 => x"58",     385 => x"78",     386 => x"96",     387 => x"B1",     388 => x"C3",     389 => x"C7",     390 => x"C2",     391 => x"B3", 
    392 => x"A2",     393 => x"8F",     394 => x"7C",     395 => x"6C",     396 => x"5C",     397 => x"51",     398 => x"48",     399 => x"48", 
    400 => x"4B",     401 => x"53",     402 => x"5F",     403 => x"6A",     404 => x"78",     405 => x"7F",     406 => x"85",     407 => x"85", 
    408 => x"87",     409 => x"8F",     410 => x"8C",     411 => x"86",     412 => x"77",     413 => x"61",     414 => x"44",     415 => x"37", 
    416 => x"2F",     417 => x"36",     418 => x"4A",     419 => x"68",     420 => x"8C",     421 => x"AC",     422 => x"C6",     423 => x"D2", 
    424 => x"D1",     425 => x"C4",     426 => x"B0",     427 => x"9B",     428 => x"82",     429 => x"6F",     430 => x"5E",     431 => x"52", 
    432 => x"4A",     433 => x"46",     434 => x"49",     435 => x"4D",     436 => x"59",     437 => x"64",     438 => x"70",     439 => x"7B", 
    440 => x"7F",     441 => x"83",     442 => x"7F",     443 => x"86",     444 => x"8B",     445 => x"87",     446 => x"7D",     447 => x"6D", 
    448 => x"52",     449 => x"3B",     450 => x"31",     451 => x"2E",     452 => x"3E",     453 => x"56",     454 => x"7D",     455 => x"A0", 
    456 => x"BF",     457 => x"D4",     458 => x"D5",     459 => x"CD",     460 => x"B6",     461 => x"A0",     462 => x"86",     463 => x"6F", 
    464 => x"60",     465 => x"52",     466 => x"4D",     467 => x"47",     468 => x"4B",     469 => x"4F",     470 => x"58",     471 => x"65", 
    472 => x"6F",     473 => x"7C",     474 => x"82",     475 => x"87",     476 => x"84",     477 => x"81",     478 => x"89",     479 => x"89", 
    480 => x"85",     481 => x"79",     482 => x"68",     483 => x"49",     484 => x"36",     485 => x"2D",     486 => x"2F",     487 => x"45", 
    488 => x"62",     489 => x"8D",     490 => x"AE",     491 => x"CE",     492 => x"DB",     493 => x"D4",     494 => x"C3",     495 => x"A4", 
    496 => x"8C",     497 => x"70",     498 => x"5E",     499 => x"53",     500 => x"4C",     501 => x"4C",     502 => x"4B",     503 => x"55", 
    504 => x"5A",     505 => x"64",     506 => x"6D",     507 => x"75",     508 => x"7E",     509 => x"81",     510 => x"85",     511 => x"80", 
    512 => x"80",     513 => x"89",     514 => x"8A",     515 => x"87",     516 => x"79",     517 => x"66",     518 => x"44",     519 => x"34", 
    520 => x"27",     521 => x"2D",     522 => x"44",     523 => x"66",     524 => x"97",     525 => x"BA",     526 => x"DD",     527 => x"E3", 
    528 => x"DA",     529 => x"BF",     530 => x"99",     531 => x"7B",     532 => x"5C",     533 => x"51",     534 => x"4A",     535 => x"4E", 
    536 => x"53",     537 => x"59",     538 => x"64",     539 => x"66",     540 => x"6E",     541 => x"71",     542 => x"76",     543 => x"7B", 
    544 => x"7C",     545 => x"7F",     546 => x"79",     547 => x"7E",     548 => x"87",     549 => x"8B",     550 => x"85",     551 => x"75", 
    552 => x"60",     553 => x"38",     554 => x"28",     555 => x"19",     556 => x"27",     557 => x"43",     558 => x"6E",     559 => x"A4", 
    560 => x"C7",     561 => x"E9",     562 => x"E7",     563 => x"D9",     564 => x"B5",     565 => x"8C",     566 => x"6D",     567 => x"51", 
    568 => x"4E",     569 => x"4D",     570 => x"5D",     571 => x"65",     572 => x"6F",     573 => x"76",     574 => x"71",     575 => x"70", 
    576 => x"67",     577 => x"69",     578 => x"68",     579 => x"6E",     580 => x"77",     581 => x"78",     582 => x"85",     583 => x"8F", 
    584 => x"97",     585 => x"8C",     586 => x"79",     587 => x"5B",     588 => x"2F",     589 => x"1E",     590 => x"11",     591 => x"28", 
    592 => x"49",     593 => x"7D",     594 => x"B2",     595 => x"D4",     596 => x"EE",     597 => x"E1",     598 => x"CB",     599 => x"9B", 
    600 => x"72",     601 => x"55",     602 => x"44",     603 => x"4F",     604 => x"5A",     605 => x"75",     606 => x"7F",     607 => x"84", 
    608 => x"7D",     609 => x"6A",     610 => x"5E",     611 => x"4F",     612 => x"54",     613 => x"5A",     614 => x"6E",     615 => x"7F", 
    616 => x"89",     617 => x"98",     618 => x"9A",     619 => x"9B",     620 => x"83",     621 => x"6D",     622 => x"4B",     623 => x"25", 
    624 => x"1D",     625 => x"1B",     626 => x"3E",     627 => x"64",     628 => x"9B",     629 => x"CB",     630 => x"E4",     631 => x"EE", 
    632 => x"CF",     633 => x"AD",     634 => x"78",     635 => x"55",     636 => x"44",     637 => x"46",     638 => x"62",     639 => x"7A", 
    640 => x"97",     641 => x"95",     642 => x"8A",     643 => x"6B",     644 => x"4B",     645 => x"38",     646 => x"32",     647 => x"49", 
    648 => x"64",     649 => x"8D",     650 => x"A6",     651 => x"AD",     652 => x"A7",     653 => x"93",     654 => x"82",     655 => x"64", 
    656 => x"50",     657 => x"40",     658 => x"2E",     659 => x"2F",     660 => x"37",     661 => x"51",     662 => x"71",     663 => x"96", 
    664 => x"BE",     665 => x"D0",     666 => x"D7",     667 => x"C4",     668 => x"A3",     669 => x"7B",     670 => x"58",     671 => x"4D", 
    672 => x"4F",     673 => x"6B",     674 => x"85",     675 => x"9B",     676 => x"99",     677 => x"84",     678 => x"65",     679 => x"43", 
    680 => x"34",     681 => x"35",     682 => x"52",     683 => x"76",     684 => x"9D",     685 => x"B4",     686 => x"AF",     687 => x"9E", 
    688 => x"82",     689 => x"6F",     690 => x"58",     691 => x"4B",     692 => x"46",     693 => x"38",     694 => x"3E",     695 => x"42", 
    696 => x"59",     697 => x"72",     698 => x"91",     699 => x"B6",     700 => x"C2",     701 => x"CD",     702 => x"B4",     703 => x"99", 
    704 => x"72",     705 => x"55",     706 => x"51",     707 => x"58",     708 => x"7A",     709 => x"8D",     710 => x"A2",     711 => x"92", 
    712 => x"73",     713 => x"4B",     714 => x"28",     715 => x"23",     716 => x"34",     717 => x"69",     718 => x"99",     719 => x"C6", 
    720 => x"D1",     721 => x"B5",     722 => x"87",     723 => x"5C",     724 => x"4B",     725 => x"4A",     726 => x"58",     727 => x"6A", 
    728 => x"64",     729 => x"55",     730 => x"43",     731 => x"39",     732 => x"47",     733 => x"66",     734 => x"A1",     735 => x"CE", 
    736 => x"EB",     737 => x"E4",     738 => x"BB",     739 => x"85",     740 => x"4D",     741 => x"3D",     742 => x"45",     743 => x"70", 
    744 => x"9A",     745 => x"B5",     746 => x"AC",     747 => x"7E",     748 => x"48",     749 => x"17",     750 => x"0E",     751 => x"25", 
    752 => x"62",     753 => x"A0",     754 => x"CD",     755 => x"D7",     756 => x"B2",     757 => x"7F",     758 => x"50",     759 => x"42", 
    760 => x"49",     761 => x"5A",     762 => x"70",     763 => x"64",     764 => x"4F",     765 => x"36",     766 => x"2C",     767 => x"41", 
    768 => x"69",     769 => x"AD",     770 => x"D5",     771 => x"EF",     772 => x"D7",     773 => x"A5",     774 => x"6D",     775 => x"3F", 
    776 => x"42",     777 => x"58",     778 => x"91",     779 => x"B2",     780 => x"BF",     781 => x"9C",     782 => x"60",     783 => x"2B", 
    784 => x"08",     785 => x"19",     786 => x"42",     787 => x"8A",     788 => x"BA",     789 => x"D2",     790 => x"C1",     791 => x"90", 
    792 => x"59",     793 => x"37",     794 => x"41",     795 => x"62",     796 => x"88",     797 => x"9B",     798 => x"8C",     799 => x"58", 
    800 => x"2C",     801 => x"12",     802 => x"29",     803 => x"60",     804 => x"AC",     805 => x"E7",     806 => x"F4",     807 => x"DB", 
    808 => x"98",     809 => x"5E",     810 => x"35",     811 => x"3D",     812 => x"65",     813 => x"99",     814 => x"C0",     815 => x"BC", 
    816 => x"97",     817 => x"55",     818 => x"21",     819 => x"0C",     820 => x"23",     821 => x"58",     822 => x"95",     823 => x"C0", 
    824 => x"C4",     825 => x"A9",     826 => x"75",     827 => x"47",     828 => x"3C",     829 => x"52",     830 => x"81",     831 => x"9B", 
    832 => x"9F",     833 => x"79",     834 => x"38",     835 => x"11",     836 => x"07",     837 => x"3A",     838 => x"7C",     839 => x"CC", 
    840 => x"F5",     841 => x"E9",     842 => x"BB",     843 => x"70",     844 => x"49",     845 => x"38",     846 => x"5E",     847 => x"8F", 
    848 => x"B9",     849 => x"C4",     850 => x"A0",     851 => x"6E",     852 => x"2E",     853 => x"18",     854 => x"1F",     855 => x"4B", 
    856 => x"80",     857 => x"A8",     858 => x"B9",     859 => x"A4",     860 => x"87",     861 => x"5F",     862 => x"4A",     863 => x"54", 
    864 => x"73",     865 => x"9A",     866 => x"A1",     867 => x"8E",     868 => x"5E",     869 => x"22",     870 => x"0D",     871 => x"17", 
    872 => x"54",     873 => x"93",     874 => x"CE",     875 => x"E3",     876 => x"CA",     877 => x"A1",     878 => x"6B",     879 => x"58", 
    880 => x"57",     881 => x"7A",     882 => x"98",     883 => x"A9",     884 => x"A3",     885 => x"80",     886 => x"5E",     887 => x"39", 
    888 => x"35",     889 => x"3F",     890 => x"5E",     891 => x"7A",     892 => x"8D",     893 => x"98",     894 => x"8D",     895 => x"85", 
    896 => x"72",     897 => x"67",     898 => x"6A",     899 => x"79",     900 => x"8E",     901 => x"8D",     902 => x"7C",     903 => x"5A", 
    904 => x"2D",     905 => x"20",     906 => x"28",     907 => x"5A",     908 => x"8F",     909 => x"BF",     910 => x"D5",     911 => x"C1", 
    912 => x"A3",     913 => x"75",     914 => x"66",     915 => x"62",     916 => x"7A",     917 => x"93",     918 => x"9E",     919 => x"9A", 
    920 => x"7E",     921 => x"65",     922 => x"47",     923 => x"41",     924 => x"45",     925 => x"59",     926 => x"71",     927 => x"84", 
    928 => x"96",     929 => x"95",     930 => x"92",     931 => x"7D",     932 => x"69",     933 => x"67",     934 => x"71",     935 => x"89", 
    936 => x"89",     937 => x"79",     938 => x"53",     939 => x"1F",     940 => x"12",     941 => x"1C",     942 => x"5A",     943 => x"95", 
    944 => x"CD",     945 => x"E1",     946 => x"C6",     947 => x"A1",     948 => x"6C",     949 => x"63",     950 => x"62",     951 => x"84", 
    952 => x"9D",     953 => x"A7",     954 => x"9C",     955 => x"77",     956 => x"5D",     957 => x"3D",     958 => x"3D",     959 => x"42", 
    960 => x"5A",     961 => x"71",     962 => x"84",     963 => x"95",     964 => x"92",     965 => x"90",     966 => x"7E",     967 => x"6C", 
    968 => x"63",     969 => x"70",     970 => x"86",     971 => x"92",     972 => x"7F",     973 => x"61",     974 => x"29",     975 => x"0F", 
    976 => x"16",     977 => x"48",     978 => x"8E",     979 => x"C4",     980 => x"E8",     981 => x"D0",     982 => x"AE",     983 => x"7A", 
    984 => x"64",     985 => x"64",     986 => x"79",     987 => x"98",     988 => x"9D",     989 => x"99",     990 => x"79",     991 => x"62", 
    992 => x"4B",     993 => x"44",     994 => x"4C",     995 => x"56",     996 => x"6B",     997 => x"75",     998 => x"87",     999 => x"8A", 
    1000 => x"8F",     1001 => x"83",     1002 => x"6F",     1003 => x"70",     1004 => x"72",     1005 => x"8B",     1006 => x"84",     1007 => x"73", 
    1008 => x"4B",     1009 => x"15",     1010 => x"0D",     1011 => x"1B",     1012 => x"63",     1013 => x"9D",     1014 => x"D7",     1015 => x"E2", 
    1016 => x"C3",     1017 => x"9B",     1018 => x"6A",     1019 => x"68",     1020 => x"6B",     1021 => x"8F",     1022 => x"9F",     1023 => x"A2", 
    1024 => x"92",     1025 => x"71",     1026 => x"60",     1027 => x"47",     1028 => x"4A",     1029 => x"4A",     1030 => x"5B",     1031 => x"6A", 
    1032 => x"7A",     1033 => x"8E",     1034 => x"91",     1035 => x"97",     1036 => x"83",     1037 => x"70",     1038 => x"66",     1039 => x"70", 
    1040 => x"88",     1041 => x"8E",     1042 => x"7B",     1043 => x"54",     1044 => x"19",     1045 => x"08",     1046 => x"16",     1047 => x"5B", 
    1048 => x"A1",     1049 => x"D9",     1050 => x"EB",     1051 => x"C5",     1052 => x"9A",     1053 => x"68",     1054 => x"62",     1055 => x"6B", 
    1056 => x"8B",     1057 => x"A2",     1058 => x"9F",     1059 => x"90",     1060 => x"6E",     1061 => x"5C",     1062 => x"48",     1063 => x"49", 
    1064 => x"4E",     1065 => x"58",     1066 => x"67",     1067 => x"72",     1068 => x"89",     1069 => x"8F",     1070 => x"96",     1071 => x"82", 
    1072 => x"6D",     1073 => x"6A",     1074 => x"71",     1075 => x"8B",     1076 => x"85",     1077 => x"72",     1078 => x"40",     1079 => x"0C", 
    1080 => x"05",     1081 => x"1D",     1082 => x"6F",     1083 => x"AD",     1084 => x"E8",     1085 => x"E5",     1086 => x"C0",     1087 => x"8F", 
    1088 => x"64",     1089 => x"66",     1090 => x"6F",     1091 => x"97",     1092 => x"A5",     1093 => x"A7",     1094 => x"8E",     1095 => x"6C", 
    1096 => x"54",     1097 => x"3D",     1098 => x"44",     1099 => x"49",     1100 => x"61",     1101 => x"6F",     1102 => x"83",     1103 => x"92", 
    1104 => x"94",     1105 => x"93",     1106 => x"7A",     1107 => x"67",     1108 => x"65",     1109 => x"76",     1110 => x"90",     1111 => x"8C", 
    1112 => x"75",     1113 => x"3D",     1114 => x"07",     1115 => x"01",     1116 => x"1F",     1117 => x"71",     1118 => x"B4",     1119 => x"EB", 
    1120 => x"E7",     1121 => x"C1",     1122 => x"8F",     1123 => x"64",     1124 => x"63",     1125 => x"6E",     1126 => x"94",     1127 => x"A3", 
    1128 => x"A2",     1129 => x"89",     1130 => x"66",     1131 => x"4F",     1132 => x"3C",     1133 => x"45",     1134 => x"4F",     1135 => x"64", 
    1136 => x"73",     1137 => x"82",     1138 => x"8E",     1139 => x"8E",     1140 => x"8A",     1141 => x"70",     1142 => x"72",     1143 => x"74", 
    1144 => x"8B",     1145 => x"8D",     1146 => x"74",     1147 => x"4F",     1148 => x"0C",     1149 => x"03",     1150 => x"0D",     1151 => x"5A", 
    1152 => x"A1",     1153 => x"DD",     1154 => x"F2",     1155 => x"CC",     1156 => x"A6",     1157 => x"6C",     1158 => x"67",     1159 => x"67", 
    1160 => x"89",     1161 => x"A2",     1162 => x"A7",     1163 => x"9E",     1164 => x"76",     1165 => x"60",     1166 => x"3E",     1167 => x"3D", 
    1168 => x"42",     1169 => x"58",     1170 => x"72",     1171 => x"83",     1172 => x"99",     1173 => x"94",     1174 => x"94",     1175 => x"78", 
    1176 => x"66",     1177 => x"67",     1178 => x"75",     1179 => x"93",     1180 => x"89",     1181 => x"75",     1182 => x"3A",     1183 => x"06", 
    1184 => x"01",     1185 => x"1C",     1186 => x"71",     1187 => x"AF",     1188 => x"EC",     1189 => x"E5",     1190 => x"C3",     1191 => x"8E", 
    1192 => x"61",     1193 => x"5F",     1194 => x"68",     1195 => x"92",     1196 => x"A1",     1197 => x"A8",     1198 => x"8E",     1199 => x"6C", 
    1200 => x"53",     1201 => x"3B",     1202 => x"41",     1203 => x"48",     1204 => x"64",     1205 => x"74",     1206 => x"89",     1207 => x"93", 
    1208 => x"91",     1209 => x"8D",     1210 => x"71",     1211 => x"6A",     1212 => x"6A",     1213 => x"7F",     1214 => x"90",     1215 => x"80", 
    1216 => x"68",     1217 => x"28",     1218 => x"0B",     1219 => x"09",     1220 => x"38",     1221 => x"85",     1222 => x"C2",     1223 => x"F2", 
    1224 => x"DB",     1225 => x"BA",     1226 => x"7C",     1227 => x"5F",     1228 => x"5A",     1229 => x"6F",     1230 => x"98",     1231 => x"A6", 
    1232 => x"AB",     1233 => x"89",     1234 => x"6B",     1235 => x"46",     1236 => x"34",     1237 => x"3B",     1238 => x"4A",     1239 => x"6C", 
    1240 => x"7E",     1241 => x"95",     1242 => x"96",     1243 => x"93",     1244 => x"84",     1245 => x"6A",     1246 => x"64",     1247 => x"6A", 
    1248 => x"83",     1249 => x"8E",     1250 => x"7E",     1251 => x"5F",     1252 => x"23",     1253 => x"0B",     1254 => x"0C",     1255 => x"41", 
    1256 => x"89",     1257 => x"C8",     1258 => x"F2",     1259 => x"DE",     1260 => x"BB",     1261 => x"7C",     1262 => x"5D",     1263 => x"53", 
    1264 => x"6A",     1265 => x"92",     1266 => x"A6",     1267 => x"AC",     1268 => x"8C",     1269 => x"6C",     1270 => x"44",     1271 => x"31", 
    1272 => x"36",     1273 => x"4A",     1274 => x"6B",     1275 => x"82",     1276 => x"9A",     1277 => x"9A",     1278 => x"95",     1279 => x"80", 
    1280 => x"66",     1281 => x"65",     1282 => x"6F",     1283 => x"8B",     1284 => x"8F",     1285 => x"7F",     1286 => x"58",     1287 => x"1B", 
    1288 => x"09",     1289 => x"0E",     1290 => x"4D",     1291 => x"8F",     1292 => x"D3",     1293 => x"F3",     1294 => x"DF",     1295 => x"B8", 
    1296 => x"77",     1297 => x"5B",     1298 => x"4E",     1299 => x"6B",     1300 => x"90",     1301 => x"A9",     1302 => x"AE",     1303 => x"8E", 
    1304 => x"6C",     1305 => x"3E",     1306 => x"2D",     1307 => x"30",     1308 => x"49",     1309 => x"6E",     1310 => x"8A",     1311 => x"A3", 
    1312 => x"A0",     1313 => x"96",     1314 => x"77",     1315 => x"5F",     1316 => x"60",     1317 => x"6E",     1318 => x"8B",     1319 => x"87", 
    1320 => x"7A",     1321 => x"49",     1322 => x"19",     1323 => x"0A",     1324 => x"17",     1325 => x"5A",     1326 => x"97",     1327 => x"DF", 
    1328 => x"F1",     1329 => x"E2",     1330 => x"B2",     1331 => x"75",     1332 => x"56",     1333 => x"49",     1334 => x"6B",     1335 => x"8D", 
    1336 => x"AC",     1337 => x"AD",     1338 => x"8F",     1339 => x"6A",     1340 => x"3A",     1341 => x"2B",     1342 => x"2B",     1343 => x"4B", 
    1344 => x"6E",     1345 => x"90",     1346 => x"A8",     1347 => x"A5",     1348 => x"98",     1349 => x"74",     1350 => x"5E",     1351 => x"5C", 
    1352 => x"6B",     1353 => x"83",     1354 => x"80",     1355 => x"77",     1356 => x"47",     1357 => x"24",     1358 => x"14",     1359 => x"25", 
    1360 => x"5F",     1361 => x"98",     1362 => x"DC",     1363 => x"ED",     1364 => x"E6",     1365 => x"B5",     1366 => x"7D",     1367 => x"59", 
    1368 => x"46",     1369 => x"60",     1370 => x"7C",     1371 => x"9E",     1372 => x"A3",     1373 => x"92",     1374 => x"74",     1375 => x"49", 
    1376 => x"37",     1377 => x"2F",     1378 => x"45",     1379 => x"61",     1380 => x"86",     1381 => x"A3",     1382 => x"AA",     1383 => x"A4", 
    1384 => x"82",     1385 => x"6C",     1386 => x"60",     1387 => x"66",     1388 => x"6F",     1389 => x"6A",     1390 => x"65",     1391 => x"3F", 
    1392 => x"2F",     1393 => x"25",     1394 => x"3D",     1395 => x"6A",     1396 => x"9D",     1397 => x"D6",     1398 => x"E5",     1399 => x"E5", 
    1400 => x"BB",     1401 => x"8E",     1402 => x"64",     1403 => x"4D",     1404 => x"58",     1405 => x"69",     1406 => x"88",     1407 => x"91", 
    1408 => x"90",     1409 => x"7C",     1410 => x"5E",     1411 => x"4B",     1412 => x"3B",     1413 => x"42",     1414 => x"52",     1415 => x"74", 
    1416 => x"92",     1417 => x"A4",     1418 => x"A9",     1419 => x"93",     1420 => x"82",     1421 => x"73",     1422 => x"6F",     1423 => x"67", 
    1424 => x"5B",     1425 => x"4F",     1426 => x"2E",     1427 => x"28",     1428 => x"27",     1429 => x"47",     1430 => x"71",     1431 => x"A5", 
    1432 => x"D7",     1433 => x"E7",     1434 => x"E9",     1435 => x"C5",     1436 => x"9D",     1437 => x"74",     1438 => x"58",     1439 => x"56", 
    1440 => x"5B",     1441 => x"6F",     1442 => x"77",     1443 => x"7F",     1444 => x"77",     1445 => x"68",     1446 => x"5D",     1447 => x"4E", 
    1448 => x"4D",     1449 => x"50",     1450 => x"65",     1451 => x"7A",     1452 => x"8D",     1453 => x"99",     1454 => x"92",     1455 => x"8F", 
    1456 => x"86",     1457 => x"7E",     1458 => x"6C",     1459 => x"57",     1460 => x"41",     1461 => x"24",     1462 => x"23",     1463 => x"2A", 
    1464 => x"4D",     1465 => x"76",     1466 => x"A8",     1467 => x"D2",     1468 => x"E3",     1469 => x"E6",     1470 => x"CA",     1471 => x"AB", 
    1472 => x"85",     1473 => x"67",     1474 => x"5B",     1475 => x"54",     1476 => x"5C",     1477 => x"61",     1478 => x"6D",     1479 => x"6E", 
    1480 => x"6C",     1481 => x"68",     1482 => x"5D",     1483 => x"5B",     1484 => x"5A",     1485 => x"65",     1486 => x"71",     1487 => x"7D", 
    1488 => x"86",     1489 => x"85",     1490 => x"8A",     1491 => x"8A",     1492 => x"84",     1493 => x"73",     1494 => x"5E",     1495 => x"44", 
    1496 => x"2D",     1497 => x"2B",     1498 => x"36",     1499 => x"55",     1500 => x"79",     1501 => x"A4",     1502 => x"C4",     1503 => x"D5", 
    1504 => x"D7",     1505 => x"C7",     1506 => x"B1",     1507 => x"95",     1508 => x"7D",     1509 => x"6D",     1510 => x"5F",     1511 => x"5B", 
    1512 => x"57",     1513 => x"5A",     1514 => x"5A",     1515 => x"5C",     1516 => x"5E",     1517 => x"5F",     1518 => x"63",     1519 => x"67", 
    1520 => x"70",     1521 => x"77",     1522 => x"7D",     1523 => x"7E",     1524 => x"7D",     1525 => x"83",     1526 => x"83",     1527 => x"7D", 
    1528 => x"6F",     1529 => x"5F",     1530 => x"49",     1531 => x"3E",     1532 => x"41",     1533 => x"4F",     1534 => x"67",     1535 => x"81", 
    1536 => x"9D",     1537 => x"AF",     1538 => x"BA",     1539 => x"BB",     1540 => x"B4",     1541 => x"A9",     1542 => x"9A",     1543 => x"8D", 
    1544 => x"7F",     1545 => x"73",     1546 => x"68",     1547 => x"60",     1548 => x"5B",     1549 => x"57",     1550 => x"58",     1551 => x"58", 
    1552 => x"5A",     1553 => x"60",     1554 => x"66",     1555 => x"6E",     1556 => x"73",     1557 => x"79",     1558 => x"79",     1559 => x"7C", 
    1560 => x"82",     1561 => x"80",     1562 => x"7A",     1563 => x"6F",     1564 => x"62",     1565 => x"55",     1566 => x"52",     1567 => x"57", 
    1568 => x"62",     1569 => x"71",     1570 => x"82",     1571 => x"90",     1572 => x"9B",     1573 => x"A2",     1574 => x"A4",     1575 => x"A1", 
    1576 => x"9D",     1577 => x"96",     1578 => x"90",     1579 => x"89",     1580 => x"80",     1581 => x"77",     1582 => x"6F",     1583 => x"66", 
    1584 => x"60",     1585 => x"5D",     1586 => x"5A",     1587 => x"58",     1588 => x"5A",     1589 => x"5D",     1590 => x"60",     1591 => x"64", 
    1592 => x"69",     1593 => x"6F",     1594 => x"78",     1595 => x"7B",     1596 => x"79",     1597 => x"74",     1598 => x"6A",     1599 => x"60", 
    1600 => x"5D",     1601 => x"61",     1602 => x"69",     1603 => x"73",     1604 => x"7F",     1605 => x"8A",     1606 => x"92",     1607 => x"98", 
    1608 => x"9A",     1609 => x"98",     1610 => x"96",     1611 => x"94",     1612 => x"93",     1613 => x"91",     1614 => x"8D",     1615 => x"85", 
    1616 => x"7D",     1617 => x"73",     1618 => x"6D",     1619 => x"69",     1620 => x"64",     1621 => x"5F",     1622 => x"5A",     1623 => x"57", 
    1624 => x"57",     1625 => x"59",     1626 => x"5D",     1627 => x"66",     1628 => x"6F",     1629 => x"72",     1630 => x"70",     1631 => x"6C", 
    1632 => x"65",     1633 => x"62",     1634 => x"64",     1635 => x"6A",     1636 => x"71",     1637 => x"7B",     1638 => x"85",     1639 => x"8C", 
    1640 => x"90",     1641 => x"93",     1642 => x"95",     1643 => x"98",     1644 => x"9A",     1645 => x"9D",     1646 => x"9C",     1647 => x"95", 
    1648 => x"8C",     1649 => x"82",     1650 => x"7A",     1651 => x"72",     1652 => x"6D",     1653 => x"66",     1654 => x"5E",     1655 => x"58", 
    1656 => x"54",     1657 => x"53",     1658 => x"53",     1659 => x"55",     1660 => x"5A",     1661 => x"62",     1662 => x"67",     1663 => x"68", 
    1664 => x"69",     1665 => x"66",     1666 => x"65",     1667 => x"68",     1668 => x"70",     1669 => x"79",     1670 => x"81",     1671 => x"88", 
    1672 => x"8C",     1673 => x"8F",     1674 => x"92",     1675 => x"97",     1676 => x"9C",     1677 => x"A0",     1678 => x"A1",     1679 => x"9E", 
    1680 => x"97",     1681 => x"8F",     1682 => x"87",     1683 => x"7F",     1684 => x"77",     1685 => x"6D",     1686 => x"64",     1687 => x"5C", 
    1688 => x"56",     1689 => x"52",     1690 => x"51",     1691 => x"4F",     1692 => x"4F",     1693 => x"54",     1694 => x"5A",     1695 => x"60", 
    1696 => x"65",     1697 => x"68",     1698 => x"6A",     1699 => x"6C",     1700 => x"70",     1701 => x"76",     1702 => x"7E",     1703 => x"84", 
    1704 => x"8A",     1705 => x"8D",     1706 => x"91",     1707 => x"95",     1708 => x"9A",     1709 => x"9D",     1710 => x"9D",     1711 => x"9C", 
    1712 => x"98",     1713 => x"92",     1714 => x"8B",     1715 => x"84",     1716 => x"7A",     1717 => x"70",     1718 => x"67",     1719 => x"5F", 
    1720 => x"57",     1721 => x"51",     1722 => x"4D",     1723 => x"4A",     1724 => x"4B",     1725 => x"50",     1726 => x"55",     1727 => x"5A", 
    1728 => x"5F",     1729 => x"64",     1730 => x"69",     1731 => x"71",     1732 => x"79",     1733 => x"81",     1734 => x"87",     1735 => x"8C", 
    1736 => x"90",     1737 => x"94",     1738 => x"98",     1739 => x"9B",     1740 => x"9D",     1741 => x"9E",     1742 => x"9C",     1743 => x"99", 
    1744 => x"94",     1745 => x"8C",     1746 => x"84",     1747 => x"7C",     1748 => x"73",     1749 => x"6A",     1750 => x"61",     1751 => x"5A", 
    1752 => x"54",     1753 => x"50",     1754 => x"4E",     1755 => x"4E",     1756 => x"50",     1757 => x"54",     1758 => x"56",     1759 => x"5B", 
    1760 => x"60",     1761 => x"65",     1762 => x"6C",     1763 => x"75",     1764 => x"7F",     1765 => x"87",     1766 => x"8D",     1767 => x"92", 
    1768 => x"95",     1769 => x"98",     1770 => x"9B",     1771 => x"9D",     1772 => x"9D",     1773 => x"9B",     1774 => x"97",     1775 => x"91", 
    1776 => x"8A",     1777 => x"83",     1778 => x"7B",     1779 => x"73",     1780 => x"6B",     1781 => x"62",     1782 => x"5B",     1783 => x"55", 
    1784 => x"51",     1785 => x"50",     1786 => x"51",     1787 => x"53",     1788 => x"56",     1789 => x"5A",     1790 => x"5E",     1791 => x"63", 
    1792 => x"69",     1793 => x"6F",     1794 => x"76",     1795 => x"7D",     1796 => x"84",     1797 => x"89",     1798 => x"8E",     1799 => x"92", 
    1800 => x"96",     1801 => x"97",     1802 => x"98",     1803 => x"98",     1804 => x"95",     1805 => x"92",     1806 => x"8D",     1807 => x"87", 
    1808 => x"80",     1809 => x"79",     1810 => x"71",     1811 => x"69",     1812 => x"62",     1813 => x"5D",     1814 => x"58",     1815 => x"56", 
    1816 => x"56",     1817 => x"58",     1818 => x"5A",     1819 => x"5D",     1820 => x"60",     1821 => x"64",     1822 => x"68",     1823 => x"6D", 
    1824 => x"73",     1825 => x"78",     1826 => x"7D",     1827 => x"81",     1828 => x"84",     1829 => x"88",     1830 => x"8C",     1831 => x"8F", 
    1832 => x"92",     1833 => x"93",     1834 => x"93",     1835 => x"91",     1836 => x"8D",     1837 => x"8A",     1838 => x"85",     1839 => x"80", 
    1840 => x"7B",     1841 => x"75",     1842 => x"70",     1843 => x"6B",     1844 => x"67",     1845 => x"63",     1846 => x"5F",     1847 => x"5D", 
    1848 => x"5B",     1849 => x"5A",     1850 => x"5C",     1851 => x"5F",     1852 => x"62",     1853 => x"66",     1854 => x"6A",     1855 => x"6E", 
    1856 => x"72",     1857 => x"76",     1858 => x"7A",     1859 => x"7E",     1860 => x"81",     1861 => x"83",     1862 => x"84",     1863 => x"85", 
    1864 => x"86",     1865 => x"88",     1866 => x"8A",     1867 => x"8B",     1868 => x"8C",     1869 => x"8B",     1870 => x"89",     1871 => x"85", 
    1872 => x"82",     1873 => x"7D",     1874 => x"79",     1875 => x"74",     1876 => x"70",     1877 => x"6C",     1878 => x"69",     1879 => x"67", 
    1880 => x"65",     1881 => x"64",     1882 => x"62",     1883 => x"61",     1884 => x"62",     1885 => x"64",     1886 => x"66",     1887 => x"6A", 
    1888 => x"6E",     1889 => x"71",     1890 => x"73",     1891 => x"75",     1892 => x"78",     1893 => x"7A",     1894 => x"7D",     1895 => x"7F", 
    1896 => x"80",     1897 => x"81",     1898 => x"82",     1899 => x"82",     1900 => x"83",     1901 => x"84",     1902 => x"85",     1903 => x"85", 
    1904 => x"85",     1905 => x"83",     1906 => x"81",     1907 => x"7F",     1908 => x"7C",     1909 => x"78",     1910 => x"75",     1911 => x"72", 
    1912 => x"6F",     1913 => x"6D",     1914 => x"6B",     1915 => x"6A",     1916 => x"69",     1917 => x"68",     1918 => x"68",     1919 => x"68", 
    1920 => x"69",     1921 => x"6B",     1922 => x"6D",     1923 => x"6F",     1924 => x"71",     1925 => x"72",     1926 => x"73",     1927 => x"74", 
    1928 => x"76",     1929 => x"78",     1930 => x"79",     1931 => x"7A",     1932 => x"7A",     1933 => x"7B",     1934 => x"7C",     1935 => x"7D", 
    1936 => x"7E",     1937 => x"80",     1938 => x"82",     1939 => x"83",     1940 => x"82",     1941 => x"82",     1942 => x"80",     1943 => x"7D", 
    1944 => x"7B",     1945 => x"7A",     1946 => x"77",     1947 => x"75",     1948 => x"74",     1949 => x"72",     1950 => x"70",     1951 => x"6F", 
    1952 => x"6E",     1953 => x"6D",     1954 => x"6C",     1955 => x"6C",     1956 => x"6C",     1957 => x"6D",     1958 => x"6D",     1959 => x"6D", 
    1960 => x"6E",     1961 => x"6F",     1962 => x"70",     1963 => x"72",     1964 => x"73",     1965 => x"75",     1966 => x"77",     1967 => x"78", 
    1968 => x"78",     1969 => x"79",     1970 => x"7A",     1971 => x"7C",     1972 => x"7E",     1973 => x"80",     1974 => x"82",     1975 => x"83", 
    1976 => x"83",     1977 => x"82",     1978 => x"82",     1979 => x"81",     1980 => x"7F",     1981 => x"7D",     1982 => x"7C",     1983 => x"79", 
    1984 => x"77",     1985 => x"75",     1986 => x"73",     1987 => x"71",     1988 => x"70",     1989 => x"6F",     1990 => x"6F",     1991 => x"6F", 
    1992 => x"6F",     1993 => x"6F",     1994 => x"6E",     1995 => x"6D",     1996 => x"6D",     1997 => x"6D",     1998 => x"6E",     1999 => x"70", 
    2000 => x"71",     2001 => x"72",     2002 => x"72",     2003 => x"73",     2004 => x"75",     2005 => x"76",     2006 => x"79",     2007 => x"7C", 
    2008 => x"7E",     2009 => x"7E",     2010 => x"7F",     2011 => x"80",     2012 => x"80",     2013 => x"7F",     2014 => x"7E",     2015 => x"7E", 
    2016 => x"7E",     2017 => x"7D",     2018 => x"7C",     2019 => x"7B",     2020 => x"7A",     2021 => x"78",     2022 => x"77",     2023 => x"76", 
    2024 => x"74",     2025 => x"73",     2026 => x"72",     2027 => x"70",     2028 => x"6F",     2029 => x"6E",     2030 => x"6D",     2031 => x"6D", 
    2032 => x"6E",     2033 => x"6F",     2034 => x"70",     2035 => x"70",     2036 => x"70",     2037 => x"71",     2038 => x"71",     2039 => x"71", 
    2040 => x"73",     2041 => x"74",     2042 => x"75",     2043 => x"77",     2044 => x"77",     2045 => x"78",     2046 => x"79",     2047 => x"79", 
    2048 => x"7A",     2049 => x"7B",     2050 => x"7C",     2051 => x"7D",     2052 => x"7E",     2053 => x"7E",     2054 => x"7E",     2055 => x"7D", 
    2056 => x"7D",     2057 => x"7D",     2058 => x"7D",     2059 => x"7C",     2060 => x"7A",     2061 => x"78",     2062 => x"76",     2063 => x"74", 
    2064 => x"72",     2065 => x"71",     2066 => x"6F",     2067 => x"6F",     2068 => x"6E",     2069 => x"6E",     2070 => x"6E",     2071 => x"6E", 
    2072 => x"6E",     2073 => x"6F",     2074 => x"70",     2075 => x"72",     2076 => x"73",     2077 => x"75",     2078 => x"75",     2079 => x"75", 
    2080 => x"75",     2081 => x"75",     2082 => x"76",     2083 => x"77",     2084 => x"78",     2085 => x"79",     2086 => x"7A",     2087 => x"7A", 
    2088 => x"7B",     2089 => x"7B",     2090 => x"7C",     2091 => x"7E",     2092 => x"7F",     2093 => x"80",     2094 => x"80",     2095 => x"80", 
    2096 => x"7F",     2097 => x"7D",     2098 => x"7B",     2099 => x"79",     2100 => x"77",     2101 => x"75",     2102 => x"74",     2103 => x"73", 
    2104 => x"71",     2105 => x"6E",     2106 => x"6D",     2107 => x"6C",     2108 => x"6C",     2109 => x"6D",     2110 => x"6E",     2111 => x"6F", 
    2112 => x"70",     2113 => x"71",     2114 => x"71",     2115 => x"71",     2116 => x"72",     2117 => x"72",     2118 => x"73",     2119 => x"74", 
    2120 => x"75",     2121 => x"76",     2122 => x"76",     2123 => x"77",     2124 => x"78",     2125 => x"7A",     2126 => x"7C",     2127 => x"7D", 
    2128 => x"7F",     2129 => x"80",     2130 => x"80",     2131 => x"80",     2132 => x"80",     2133 => x"7F",     2134 => x"7E",     2135 => x"7D", 
    2136 => x"7C",     2137 => x"7B",     2138 => x"79",     2139 => x"77",     2140 => x"74",     2141 => x"72",     2142 => x"70",     2143 => x"6F", 
    2144 => x"6E",     2145 => x"6E",     2146 => x"6E",     2147 => x"6F",     2148 => x"6F",     2149 => x"6F",     2150 => x"6F",     2151 => x"70", 
    2152 => x"70",     2153 => x"72",     2154 => x"72",     2155 => x"73",     2156 => x"73",     2157 => x"73",     2158 => x"74",     2159 => x"75", 
    2160 => x"76",     2161 => x"77",     2162 => x"78",     2163 => x"7A",     2164 => x"7B",     2165 => x"7C",     2166 => x"7D",     2167 => x"7D", 
    2168 => x"7E",     2169 => x"7E",     2170 => x"7E",     2171 => x"7E",     2172 => x"7E",     2173 => x"7D",     2174 => x"7B",     2175 => x"7A", 
    2176 => x"78",     2177 => x"76",     2178 => x"74",     2179 => x"73",     2180 => x"72",     2181 => x"71",     2182 => x"71",     2183 => x"71", 
    2184 => x"71",     2185 => x"70",     2186 => x"70",     2187 => x"70",     2188 => x"70",     2189 => x"70",     2190 => x"71",     2191 => x"72", 
    2192 => x"73",     2193 => x"73",     2194 => x"72",     2195 => x"73",     2196 => x"74",     2197 => x"75",     2198 => x"76",     2199 => x"78", 
    2200 => x"78",     2201 => x"78",     2202 => x"78",     2203 => x"78",     2204 => x"7A",     2205 => x"7B",     2206 => x"7C",     2207 => x"7D", 
    2208 => x"7E",     2209 => x"7F",     2210 => x"7E",     2211 => x"7E",     2212 => x"7D",     2213 => x"7C",     2214 => x"7A",     2215 => x"79", 
    2216 => x"77",     2217 => x"76",     2218 => x"74",     2219 => x"73",     2220 => x"72",     2221 => x"71",     2222 => x"71",     2223 => x"70", 
    2224 => x"71",     2225 => x"71",     2226 => x"71",     2227 => x"72",     2228 => x"72",     2229 => x"72",     2230 => x"73",     2231 => x"73", 
    2232 => x"73",     2233 => x"74",     2234 => x"74",     2235 => x"74",     2236 => x"73",     2237 => x"73",     2238 => x"73",     2239 => x"74", 
    2240 => x"75",     2241 => x"76",     2242 => x"78",     2243 => x"7A",     2244 => x"7B",     2245 => x"7C",     2246 => x"7D",     2247 => x"7D", 
    2248 => x"7E",     2249 => x"7E",     2250 => x"7E",     2251 => x"7E",     2252 => x"7C",     2253 => x"7B",     2254 => x"79",     2255 => x"78", 
    2256 => x"76",     2257 => x"75",     2258 => x"74",     2259 => x"74",     2260 => x"73",     2261 => x"72",     2262 => x"72",     2263 => x"72", 
    2264 => x"71",     2265 => x"71",     2266 => x"71",     2267 => x"72",     2268 => x"73",     2269 => x"74",     2270 => x"74",     2271 => x"74", 
    2272 => x"74",     2273 => x"75",     2274 => x"75",     2275 => x"75",     2276 => x"75",     2277 => x"76",     2278 => x"76",     2279 => x"76", 
    2280 => x"78",     2281 => x"78",     2282 => x"77",     2283 => x"78",     2284 => x"7A",     2285 => x"7B",     2286 => x"7C",     2287 => x"7C", 
    2288 => x"7C",     2289 => x"7C",     2290 => x"7B",     2291 => x"7B",     2292 => x"7A",     2293 => x"79",     2294 => x"78",     2295 => x"76", 
    2296 => x"75",     2297 => x"73",     2298 => x"72",     2299 => x"72",     2300 => x"71",     2301 => x"72",     2302 => x"72",     2303 => x"72", 
    2304 => x"72",     2305 => x"73",     2306 => x"73",     2307 => x"73",     2308 => x"73",     2309 => x"74",     2310 => x"75",     2311 => x"74", 
    2312 => x"74",     2313 => x"74",     2314 => x"74",     2315 => x"74",     2316 => x"73",     2317 => x"73",     2318 => x"74",     2319 => x"75", 
    2320 => x"77",     2321 => x"78",     2322 => x"79",     2323 => x"7A",     2324 => x"7A",     2325 => x"7A",     2326 => x"7A",     2327 => x"79", 
    2328 => x"7B",     2329 => x"7B",     2330 => x"7C",     2331 => x"7C",     2332 => x"7B",     2333 => x"7A",     2334 => x"79",     2335 => x"79", 
    2336 => x"77",     2337 => x"76",     2338 => x"74",     2339 => x"73",     2340 => x"72",     2341 => x"72",     2342 => x"72",     2343 => x"73", 
    2344 => x"72",     2345 => x"72",     2346 => x"72",     2347 => x"72",     2348 => x"73",     2349 => x"74",     2350 => x"76",     2351 => x"76", 
    2352 => x"75",     2353 => x"75",     2354 => x"76",     2355 => x"76",     2356 => x"76",     2357 => x"75",     2358 => x"74",     2359 => x"75", 
    2360 => x"75",     2361 => x"77",     2362 => x"77",     2363 => x"77",     2364 => x"77",     2365 => x"77",     2366 => x"77",     2367 => x"77", 
    2368 => x"78",     2369 => x"79",     2370 => x"7A",     2371 => x"79",     2372 => x"7A",     2373 => x"79",     2374 => x"7A",     2375 => x"7B", 
    2376 => x"7A",     2377 => x"7A",     2378 => x"79",     2379 => x"78",     2380 => x"75",     2381 => x"74",     2382 => x"73",     2383 => x"73", 
    2384 => x"73",     2385 => x"74",     2386 => x"75",     2387 => x"75",     2388 => x"75",     2389 => x"74",     2390 => x"74",     2391 => x"74", 
    2392 => x"75",     2393 => x"76",     2394 => x"76",     2395 => x"77",     2396 => x"77",     2397 => x"76",     2398 => x"76",     2399 => x"74", 
    2400 => x"73",     2401 => x"74",     2402 => x"75",     2403 => x"76",     2404 => x"77",     2405 => x"76",     2406 => x"76",     2407 => x"76", 
    2408 => x"76",     2409 => x"76",     2410 => x"76",     2411 => x"78",     2412 => x"79",     2413 => x"7A",     2414 => x"7A",     2415 => x"7B", 
    2416 => x"7A",     2417 => x"7C",     2418 => x"7D",     2419 => x"7C",     2420 => x"7A",     2421 => x"78",     2422 => x"77",     2423 => x"75", 
    2424 => x"74",     2425 => x"73",     2426 => x"73",     2427 => x"73",     2428 => x"74",     2429 => x"74",     2430 => x"73",     2431 => x"74", 
    2432 => x"73",     2433 => x"73",     2434 => x"73",     2435 => x"72",     2436 => x"71",     2437 => x"71",     2438 => x"71",     2439 => x"72", 
    2440 => x"73",     2441 => x"74",     2442 => x"75",     2443 => x"74",     2444 => x"74",     2445 => x"73",     2446 => x"73",     2447 => x"74", 
    2448 => x"74",     2449 => x"75",     2450 => x"76",     2451 => x"79",     2452 => x"79",     2453 => x"7B",     2454 => x"7C",     2455 => x"7E", 
    2456 => x"7E",     2457 => x"7E",     2458 => x"7D",     2459 => x"7B",     2460 => x"7A",     2461 => x"7A",     2462 => x"7A",     2463 => x"7A", 
    2464 => x"7A",     2465 => x"79",     2466 => x"77",     2467 => x"75",     2468 => x"73",     2469 => x"73",     2470 => x"73",     2471 => x"74", 
    2472 => x"74",     2473 => x"74",     2474 => x"73",     2475 => x"73",     2476 => x"73",     2477 => x"72",     2478 => x"70",     2479 => x"6F", 
    2480 => x"6E",     2481 => x"6E",     2482 => x"6F",     2483 => x"70",     2484 => x"70",     2485 => x"71",     2486 => x"73",     2487 => x"74", 
    2488 => x"74",     2489 => x"75",     2490 => x"76",     2491 => x"78",     2492 => x"79",     2493 => x"7B",     2494 => x"7C",     2495 => x"7D", 
    2496 => x"7D",     2497 => x"7D",     2498 => x"7E",     2499 => x"7F",     2500 => x"80",     2501 => x"80",     2502 => x"7F",     2503 => x"7E", 
    2504 => x"7C",     2505 => x"79",     2506 => x"76",     2507 => x"74",     2508 => x"73",     2509 => x"74",     2510 => x"74",     2511 => x"74", 
    2512 => x"73",     2513 => x"72",     2514 => x"71",     2515 => x"70",     2516 => x"70",     2517 => x"6F",     2518 => x"6E",     2519 => x"6E", 
    2520 => x"6E",     2521 => x"6F",     2522 => x"70",     2523 => x"70",     2524 => x"71",     2525 => x"72",     2526 => x"74",     2527 => x"75", 
    2528 => x"77",     2529 => x"78",     2530 => x"7A",     2531 => x"7C",     2532 => x"7E",     2533 => x"80",     2534 => x"81",     2535 => x"81", 
    2536 => x"82",     2537 => x"83",     2538 => x"84",     2539 => x"84",     2540 => x"82",     2541 => x"80",     2542 => x"7D",     2543 => x"7A", 
    2544 => x"78",     2545 => x"75",     2546 => x"72",     2547 => x"70",     2548 => x"6F",     2549 => x"6E",     2550 => x"6E",     2551 => x"6E", 
    2552 => x"6D",     2553 => x"6B",     2554 => x"6A",     2555 => x"6A",     2556 => x"6A",     2557 => x"6B",     2558 => x"6C",     2559 => x"6D", 
    2560 => x"6F",     2561 => x"71",     2562 => x"72",     2563 => x"72",     2564 => x"73",     2565 => x"73",     2566 => x"75",     2567 => x"77", 
    2568 => x"7B",     2569 => x"7F",     2570 => x"82",     2571 => x"84",     2572 => x"84",     2573 => x"85",     2574 => x"84",     2575 => x"84", 
    2576 => x"83",     2577 => x"83",     2578 => x"82",     2579 => x"7F",     2580 => x"7C",     2581 => x"77",     2582 => x"72",     2583 => x"6D", 
    2584 => x"69",     2585 => x"67",     2586 => x"68",     2587 => x"68",     2588 => x"69",     2589 => x"6A",     2590 => x"69",     2591 => x"6B", 
    2592 => x"6B",     2593 => x"6E",     2594 => x"70",     2595 => x"73",     2596 => x"76",     2597 => x"78",     2598 => x"79",     2599 => x"7A", 
    2600 => x"7B",     2601 => x"7C",     2602 => x"7D",     2603 => x"7F",     2604 => x"81",     2605 => x"85",     2606 => x"88",     2607 => x"8C", 
    2608 => x"8E",     2609 => x"90",     2610 => x"8F",     2611 => x"8E",     2612 => x"8A",     2613 => x"85",     2614 => x"7F",     2615 => x"78", 
    2616 => x"71",     2617 => x"6B",     2618 => x"65",     2619 => x"62",     2620 => x"60",     2621 => x"60",     2622 => x"60",     2623 => x"60", 
    2624 => x"5F",     2625 => x"60",     2626 => x"63",     2627 => x"66",     2628 => x"6A",     2629 => x"6C",     2630 => x"6E",     2631 => x"6D", 
    2632 => x"6C",     2633 => x"69",     2634 => x"66",     2635 => x"64",     2636 => x"65",     2637 => x"69",     2638 => x"70",     2639 => x"7B", 
    2640 => x"87",     2641 => x"92",     2642 => x"98",     2643 => x"98",     2644 => x"95",     2645 => x"8E",     2646 => x"85",     2647 => x"7C", 
    2648 => x"73",     2649 => x"6B",     2650 => x"64",     2651 => x"60",     2652 => x"5D",     2653 => x"5B",     2654 => x"5A",     2655 => x"5A", 
    2656 => x"5D",     2657 => x"62",     2658 => x"69",     2659 => x"71",     2660 => x"7A",     2661 => x"80",     2662 => x"84",     2663 => x"84", 
    2664 => x"81",     2665 => x"7A",     2666 => x"73",     2667 => x"6E",     2668 => x"6E",     2669 => x"76",     2670 => x"85",     2671 => x"95", 
    2672 => x"A6",     2673 => x"B1",     2674 => x"B6",     2675 => x"B4",     2676 => x"AA",     2677 => x"9B",     2678 => x"8A",     2679 => x"79", 
    2680 => x"6B",     2681 => x"5F",     2682 => x"56",     2683 => x"50",     2684 => x"4D",     2685 => x"4D",     2686 => x"50",     2687 => x"55", 
    2688 => x"5C",     2689 => x"65",     2690 => x"70",     2691 => x"7B",     2692 => x"83",     2693 => x"84",     2694 => x"7E",     2695 => x"73", 
    2696 => x"67",     2697 => x"61",     2698 => x"62",     2699 => x"6F",     2700 => x"83",     2701 => x"9B",     2702 => x"B2",     2703 => x"C1", 
    2704 => x"C8",     2705 => x"C4",     2706 => x"B8",     2707 => x"A6",     2708 => x"91",     2709 => x"7D",     2710 => x"6C",     2711 => x"60", 
    2712 => x"57",     2713 => x"52",     2714 => x"4F",     2715 => x"4F",     2716 => x"52",     2717 => x"56",     2718 => x"5F",     2719 => x"6B", 
    2720 => x"78",     2721 => x"81",     2722 => x"85",     2723 => x"81",     2724 => x"74",     2725 => x"67",     2726 => x"5B",     2727 => x"57", 
    2728 => x"5F",     2729 => x"71",     2730 => x"87",     2731 => x"9C",     2732 => x"AD",     2733 => x"B5",     2734 => x"B3",     2735 => x"A9", 
    2736 => x"97",     2737 => x"82",     2738 => x"6B",     2739 => x"56",     2740 => x"46",     2741 => x"3C",     2742 => x"37",     2743 => x"36", 
    2744 => x"39",     2745 => x"3B",     2746 => x"43",     2747 => x"50",     2748 => x"61",     2749 => x"72",     2750 => x"7C",     2751 => x"81", 
    2752 => x"79",     2753 => x"6E",     2754 => x"64",     2755 => x"5D",     2756 => x"61",     2757 => x"6F",     2758 => x"85",     2759 => x"9F", 
    2760 => x"B7",     2761 => x"C8",     2762 => x"CE",     2763 => x"CA",     2764 => x"BB",     2765 => x"A7",     2766 => x"8E",     2767 => x"76", 
    2768 => x"60",     2769 => x"50",     2770 => x"47",     2771 => x"43",     2772 => x"43",     2773 => x"45",     2774 => x"48",     2775 => x"50", 
    2776 => x"5C",     2777 => x"6A",     2778 => x"75",     2779 => x"79",     2780 => x"75",     2781 => x"67",     2782 => x"5A",     2783 => x"4F", 
    2784 => x"4D",     2785 => x"58",     2786 => x"6C",     2787 => x"86",     2788 => x"A0",     2789 => x"B6",     2790 => x"C2",     2791 => x"C2", 
    2792 => x"B8",     2793 => x"A5",     2794 => x"8F",     2795 => x"76",     2796 => x"5F",     2797 => x"4C",     2798 => x"3F",     2799 => x"38", 
    2800 => x"36",     2801 => x"38",     2802 => x"3B",     2803 => x"3D",     2804 => x"46",     2805 => x"55",     2806 => x"64",     2807 => x"71", 
    2808 => x"77",     2809 => x"73",     2810 => x"63",     2811 => x"54",     2812 => x"49",     2813 => x"47",     2814 => x"56",     2815 => x"6F", 
    2816 => x"8F",     2817 => x"AD",     2818 => x"C7",     2819 => x"D5",     2820 => x"D4",     2821 => x"CB",     2822 => x"B7",     2823 => x"A1", 
    2824 => x"89",     2825 => x"74",     2826 => x"63",     2827 => x"57",     2828 => x"51",     2829 => x"4F",     2830 => x"53",     2831 => x"56", 
    2832 => x"59",     2833 => x"5C",     2834 => x"65",     2835 => x"72",     2836 => x"7D",     2837 => x"85",     2838 => x"83",     2839 => x"78", 
    2840 => x"64",     2841 => x"53",     2842 => x"48",     2843 => x"4B",     2844 => x"5F",     2845 => x"7D",     2846 => x"A1",     2847 => x"C1", 
    2848 => x"D8",     2849 => x"DF",     2850 => x"D7",     2851 => x"C5",     2852 => x"AB",     2853 => x"91",     2854 => x"78",     2855 => x"66", 
    2856 => x"5A",     2857 => x"53",     2858 => x"53",     2859 => x"55",     2860 => x"5C",     2861 => x"60",     2862 => x"62",     2863 => x"62", 
    2864 => x"67",     2865 => x"73",     2866 => x"7F",     2867 => x"8A",     2868 => x"8A",     2869 => x"84",     2870 => x"6E",     2871 => x"5C", 
    2872 => x"4E",     2873 => x"4A",     2874 => x"5C",     2875 => x"78",     2876 => x"A2",     2877 => x"C6",     2878 => x"E5",     2879 => x"F1", 
    2880 => x"E6",     2881 => x"D1",     2882 => x"AE",     2883 => x"8F",     2884 => x"71",     2885 => x"5D",     2886 => x"52",     2887 => x"4D", 
    2888 => x"52",     2889 => x"54",     2890 => x"5B",     2891 => x"5D",     2892 => x"5E",     2893 => x"5A",     2894 => x"52",     2895 => x"57", 
    2896 => x"5E",     2897 => x"6B",     2898 => x"74",     2899 => x"75",     2900 => x"6C",     2901 => x"50",     2902 => x"40",     2903 => x"2B", 
    2904 => x"2A",     2905 => x"3D",     2906 => x"5F",     2907 => x"8F",     2908 => x"B7",     2909 => x"DC",     2910 => x"E2",     2911 => x"D3", 
    2912 => x"B5",     2913 => x"89",     2914 => x"65",     2915 => x"47",     2916 => x"3C",     2917 => x"3B",     2918 => x"43",     2919 => x"52", 
    2920 => x"5A",     2921 => x"63",     2922 => x"63",     2923 => x"61",     2924 => x"5A",     2925 => x"51",     2926 => x"57",     2927 => x"62", 
    2928 => x"75",     2929 => x"83",     2930 => x"87",     2931 => x"81",     2932 => x"61",     2933 => x"4B",     2934 => x"33",     2935 => x"2D", 
    2936 => x"41",     2937 => x"65",     2938 => x"9B",     2939 => x"C7",     2940 => x"F1",     2941 => x"FD",     2942 => x"EE",     2943 => x"CD", 
    2944 => x"9A",     2945 => x"71",     2946 => x"4E",     2947 => x"43",     2948 => x"46",     2949 => x"54",     2950 => x"69",     2951 => x"74", 
    2952 => x"7F",     2953 => x"7C",     2954 => x"75",     2955 => x"6B",     2956 => x"5D",     2957 => x"57",     2958 => x"5F",     2959 => x"72", 
    2960 => x"85",     2961 => x"90",     2962 => x"8F",     2963 => x"79",     2964 => x"54",     2965 => x"39",     2966 => x"22",     2967 => x"26", 
    2968 => x"42",     2969 => x"73",     2970 => x"A9",     2971 => x"D8",     2972 => x"F9",     2973 => x"F6",     2974 => x"DA",     2975 => x"A8", 
    2976 => x"6F",     2977 => x"41",     2978 => x"23",     2979 => x"23",     2980 => x"32",     2981 => x"4E",     2982 => x"68",     2983 => x"7A", 
    2984 => x"82",     2985 => x"78",     2986 => x"6B",     2987 => x"59",     2988 => x"49",     2989 => x"40",     2990 => x"4A",     2991 => x"61", 
    2992 => x"77",     2993 => x"8A",     2994 => x"8A",     2995 => x"7B",     2996 => x"54",     2997 => x"37",     2998 => x"1E",     2999 => x"1D", 
    3000 => x"3B",     3001 => x"68",     3002 => x"A2",     3003 => x"D0",     3004 => x"F4",     3005 => x"F9",     3006 => x"E1",     3007 => x"B8", 
    3008 => x"7E",     3009 => x"50",     3010 => x"30",     3011 => x"2D",     3012 => x"40",     3013 => x"5E",     3014 => x"80",     3015 => x"93", 
    3016 => x"9B",     3017 => x"92",     3018 => x"7F",     3019 => x"6B",     3020 => x"59",     3021 => x"52",     3022 => x"52",     3023 => x"69", 
    3024 => x"84",     3025 => x"9C",     3026 => x"A8",     3027 => x"9C",     3028 => x"83",     3029 => x"55",     3030 => x"39",     3031 => x"26", 
    3032 => x"2E",     3033 => x"52",     3034 => x"80",     3035 => x"B9",     3036 => x"DD",     3037 => x"F5",     3038 => x"EF",     3039 => x"D0", 
    3040 => x"A5",     3041 => x"6F",     3042 => x"4B",     3043 => x"32",     3044 => x"36",     3045 => x"4C",     3046 => x"68",     3047 => x"88", 
    3048 => x"95",     3049 => x"99",     3050 => x"88",     3051 => x"72",     3052 => x"5D",     3053 => x"4D",     3054 => x"4F",     3055 => x"54", 
    3056 => x"6A",     3057 => x"85",     3058 => x"99",     3059 => x"A5",     3060 => x"96",     3061 => x"82",     3062 => x"55",     3063 => x"34", 
    3064 => x"24",     3065 => x"23",     3066 => x"47",     3067 => x"70",     3068 => x"AC",     3069 => x"D5",     3070 => x"EE",     3071 => x"F0", 
    3072 => x"CD",     3073 => x"A6",     3074 => x"71",     3075 => x"4C",     3076 => x"32",     3077 => x"2E",     3078 => x"43",     3079 => x"59", 
    3080 => x"79",     3081 => x"89",     3082 => x"8F",     3083 => x"84",     3084 => x"6E",     3085 => x"5F",     3086 => x"4E",     3087 => x"50", 
    3088 => x"58",     3089 => x"67",     3090 => x"7A",     3091 => x"8D",     3092 => x"9B",     3093 => x"99",     3094 => x"88",     3095 => x"6E", 
    3096 => x"4B",     3097 => x"2C",     3098 => x"24",     3099 => x"2B",     3100 => x"4B",     3101 => x"76",     3102 => x"AA",     3103 => x"D0", 
    3104 => x"E1",     3105 => x"E0",     3106 => x"C2",     3107 => x"9B",     3108 => x"6D",     3109 => x"4B",     3110 => x"38",     3111 => x"34", 
    3112 => x"47",     3113 => x"5E",     3114 => x"7A",     3115 => x"8B",     3116 => x"8F",     3117 => x"86",     3118 => x"71",     3119 => x"61", 
    3120 => x"56",     3121 => x"59",     3122 => x"65",     3123 => x"77",     3124 => x"86",     3125 => x"8E",     3126 => x"96",     3127 => x"8F", 
    3128 => x"83",     3129 => x"6A",     3130 => x"54",     3131 => x"3A",     3132 => x"2C",     3133 => x"35",     3134 => x"47",     3135 => x"6F", 
    3136 => x"96",     3137 => x"C0",     3138 => x"D6",     3139 => x"DA",     3140 => x"CF",     3141 => x"AA",     3142 => x"88",     3143 => x"60", 
    3144 => x"48",     3145 => x"3E",     3146 => x"42",     3147 => x"5A",     3148 => x"6E",     3149 => x"86",     3150 => x"8E",     3151 => x"8C", 
    3152 => x"7F",     3153 => x"6A",     3154 => x"5E",     3155 => x"54",     3156 => x"5C",     3157 => x"6A",     3158 => x"7C",     3159 => x"8A", 
    3160 => x"94",     3161 => x"98",     3162 => x"8E",     3163 => x"79",     3164 => x"5D",     3165 => x"40",     3166 => x"22",     3167 => x"1F", 
    3168 => x"2A",     3169 => x"4D",     3170 => x"7D",     3171 => x"B1",     3172 => x"DE",     3173 => x"ED",     3174 => x"EB",     3175 => x"CA", 
    3176 => x"9D",     3177 => x"70",     3178 => x"49",     3179 => x"3A",     3180 => x"37",     3181 => x"4B",     3182 => x"65",     3183 => x"7F", 
    3184 => x"8F",     3185 => x"8D",     3186 => x"83",     3187 => x"69",     3188 => x"57",     3189 => x"4D",     3190 => x"51",     3191 => x"64", 
    3192 => x"7A",     3193 => x"8E",     3194 => x"93",     3195 => x"98",     3196 => x"8E",     3197 => x"7E",     3198 => x"62",     3199 => x"49", 
    3200 => x"2F",     3201 => x"16",     3202 => x"21",     3203 => x"31",     3204 => x"61",     3205 => x"94",     3206 => x"CC",     3207 => x"F5", 
    3208 => x"FA",     3209 => x"F1",     3210 => x"BF",     3211 => x"8C",     3212 => x"59",     3213 => x"37",     3214 => x"2F",     3215 => x"35", 
    3216 => x"57",     3217 => x"71",     3218 => x"8C",     3219 => x"95",     3220 => x"8C",     3221 => x"7B",     3222 => x"5D",     3223 => x"52", 
    3224 => x"4C",     3225 => x"5A",     3226 => x"71",     3227 => x"85",     3228 => x"93",     3229 => x"90",     3230 => x"92",     3231 => x"84", 
    3232 => x"77",     3233 => x"5F",     3234 => x"4B",     3235 => x"34",     3236 => x"23",     3237 => x"30",     3238 => x"40",     3239 => x"6F", 
    3240 => x"9C",     3241 => x"D0",     3242 => x"F1",     3243 => x"F4",     3244 => x"E7",     3245 => x"B1",     3246 => x"81",     3247 => x"4E", 
    3248 => x"34",     3249 => x"33",     3250 => x"41",     3251 => x"68",     3252 => x"7F",     3253 => x"96",     3254 => x"94",     3255 => x"86", 
    3256 => x"70",     3257 => x"54",     3258 => x"4F",     3259 => x"50",     3260 => x"68",     3261 => x"82",     3262 => x"97",     3263 => x"9D", 
    3264 => x"90",     3265 => x"8B",     3266 => x"78",     3267 => x"70",     3268 => x"5C",     3269 => x"50",     3270 => x"3C",     3271 => x"27", 
    3272 => x"30",     3273 => x"38",     3274 => x"65",     3275 => x"91",     3276 => x"CA",     3277 => x"F1",     3278 => x"F5",     3279 => x"EB", 
    3280 => x"B3",     3281 => x"82",     3282 => x"4B",     3283 => x"33",     3284 => x"35",     3285 => x"44",     3286 => x"70",     3287 => x"87", 
    3288 => x"9C",     3289 => x"93",     3290 => x"7E",     3291 => x"66",     3292 => x"48",     3293 => x"49",     3294 => x"4F",     3295 => x"6E", 
    3296 => x"89",     3297 => x"9B",     3298 => x"9D",     3299 => x"83",     3300 => x"7A",     3301 => x"66",     3302 => x"65",     3303 => x"5D", 
    3304 => x"56",     3305 => x"4F",     3306 => x"30",     3307 => x"32",     3308 => x"2E",     3309 => x"51",     3310 => x"7F",     3311 => x"B6", 
    3312 => x"F1",     3313 => x"FB",     3314 => x"FC",     3315 => x"C7",     3316 => x"8B",     3317 => x"50",     3318 => x"29",     3319 => x"2F", 
    3320 => x"3E",     3321 => x"71",     3322 => x"91",     3323 => x"A4",     3324 => x"9D",     3325 => x"7A",     3326 => x"5F",     3327 => x"39", 
    3328 => x"38",     3329 => x"44",     3330 => x"65",     3331 => x"8B",     3332 => x"9F",     3333 => x"A7",     3334 => x"88",     3335 => x"73", 
    3336 => x"61",     3337 => x"5C",     3338 => x"64",     3339 => x"60",     3340 => x"66",     3341 => x"45",     3342 => x"3A",     3343 => x"31", 
    3344 => x"3C",     3345 => x"6A",     3346 => x"9B",     3347 => x"E3",     3348 => x"FA",     3349 => x"FF",     3350 => x"D8",     3351 => x"94", 
    3352 => x"5A",     3353 => x"27",     3354 => x"2B",     3355 => x"3E",     3356 => x"6F",     3357 => x"99",     3358 => x"A7",     3359 => x"A0", 
    3360 => x"74",     3361 => x"50",     3362 => x"2B",     3363 => x"28",     3364 => x"41",     3365 => x"68",     3366 => x"98",     3367 => x"AF", 
    3368 => x"B7",     3369 => x"99",     3370 => x"73",     3371 => x"5F",     3372 => x"53",     3373 => x"63",     3374 => x"68",     3375 => x"73", 
    3376 => x"63",     3377 => x"3F",     3378 => x"32",     3379 => x"23",     3380 => x"47",     3381 => x"76",     3382 => x"BD",     3383 => x"F3", 
    3384 => x"FD",     3385 => x"F1",     3386 => x"AE",     3387 => x"72",     3388 => x"38",     3389 => x"26",     3390 => x"3D",     3391 => x"61", 
    3392 => x"99",     3393 => x"AC",     3394 => x"AA",     3395 => x"80",     3396 => x"4E",     3397 => x"2F",     3398 => x"20",     3399 => x"40", 
    3400 => x"69",     3401 => x"9F",     3402 => x"BD",     3403 => x"BF",     3404 => x"A8",     3405 => x"72",     3406 => x"54",     3407 => x"47", 
    3408 => x"56",     3409 => x"70",     3410 => x"7B",     3411 => x"7F",     3412 => x"54",     3413 => x"33",     3414 => x"1C",     3415 => x"21", 
    3416 => x"55",     3417 => x"91",     3418 => x"E0",     3419 => x"FD",     3420 => x"FD",     3421 => x"CF",     3422 => x"85",     3423 => x"4D", 
    3424 => x"23",     3425 => x"36",     3426 => x"58",     3427 => x"8E",     3428 => x"B3",     3429 => x"B0",     3430 => x"97",     3431 => x"5C", 
    3432 => x"37",     3433 => x"21",     3434 => x"31",     3435 => x"5F",     3436 => x"8E",     3437 => x"B8",     3438 => x"BA",     3439 => x"AA", 
    3440 => x"7D",     3441 => x"50",     3442 => x"43",     3443 => x"4B",     3444 => x"6F",     3445 => x"86",     3446 => x"8D",     3447 => x"79", 
    3448 => x"45",     3449 => x"28",     3450 => x"15",     3451 => x"35",     3452 => x"6E",     3453 => x"B4",     3454 => x"F4",     3455 => x"FC", 
    3456 => x"ED",     3457 => x"AB",     3458 => x"6C",     3459 => x"3B",     3460 => x"2C",     3461 => x"4C",     3462 => x"72",     3463 => x"A4", 
    3464 => x"B0",     3465 => x"A2",     3466 => x"77",     3467 => x"42",     3468 => x"2A",     3469 => x"25",     3470 => x"49",     3471 => x"76", 
    3472 => x"A1",     3473 => x"B8",     3474 => x"AC",     3475 => x"93",     3476 => x"63",     3477 => x"46",     3478 => x"45",     3479 => x"5E", 
    3480 => x"85",     3481 => x"95",     3482 => x"91",     3483 => x"6B",     3484 => x"33",     3485 => x"18",     3486 => x"14",     3487 => x"45", 
    3488 => x"86",     3489 => x"CF",     3490 => x"FE",     3491 => x"F6",     3492 => x"D3",     3493 => x"8A",     3494 => x"54",     3495 => x"31", 
    3496 => x"39",     3497 => x"62",     3498 => x"88",     3499 => x"AB",     3500 => x"A5",     3501 => x"89",     3502 => x"5A",     3503 => x"34", 
    3504 => x"2C",     3505 => x"39",     3506 => x"64",     3507 => x"8D",     3508 => x"AD",     3509 => x"B1",     3510 => x"9C",     3511 => x"80", 
    3512 => x"59",     3513 => x"48",     3514 => x"53",     3515 => x"70",     3516 => x"91",     3517 => x"96",     3518 => x"87",     3519 => x"5B", 
    3520 => x"29",     3521 => x"18",     3522 => x"20",     3523 => x"58",     3524 => x"97",     3525 => x"D7",     3526 => x"F5",     3527 => x"E3", 
    3528 => x"BA",     3529 => x"78",     3530 => x"4E",     3531 => x"38",     3532 => x"4B",     3533 => x"72",     3534 => x"92",     3535 => x"A7", 
    3536 => x"96",     3537 => x"78",     3538 => x"4D",     3539 => x"34",     3540 => x"37",     3541 => x"4B",     3542 => x"74",     3543 => x"93", 
    3544 => x"A7",     3545 => x"A3",     3546 => x"8F",     3547 => x"76",     3548 => x"58",     3549 => x"50",     3550 => x"5D",     3551 => x"76", 
    3552 => x"8E",     3553 => x"8C",     3554 => x"79",     3555 => x"4F",     3556 => x"26",     3557 => x"1D",     3558 => x"2D",     3559 => x"65", 
    3560 => x"9E",     3561 => x"D7",     3562 => x"EC",     3563 => x"D7",     3564 => x"B0",     3565 => x"76",     3566 => x"55",     3567 => x"46", 
    3568 => x"5A",     3569 => x"7A",     3570 => x"91",     3571 => x"9F",     3572 => x"8C",     3573 => x"73",     3574 => x"51",     3575 => x"40", 
    3576 => x"45",     3577 => x"55",     3578 => x"77",     3579 => x"8E",     3580 => x"9E",     3581 => x"98",     3582 => x"87",     3583 => x"73", 
    3584 => x"5B",     3585 => x"56",     3586 => x"63",     3587 => x"7B",     3588 => x"8E",     3589 => x"88",     3590 => x"71",     3591 => x"46", 
    3592 => x"1F",     3593 => x"1C",     3594 => x"33",     3595 => x"6F",     3596 => x"AA",     3597 => x"DF",     3598 => x"F0",     3599 => x"D8", 
    3600 => x"AF",     3601 => x"77",     3602 => x"56",     3603 => x"4A",     3604 => x"5E",     3605 => x"7E",     3606 => x"91",     3607 => x"9A", 
    3608 => x"84",     3609 => x"69",     3610 => x"4A",     3611 => x"3C",     3612 => x"46",     3613 => x"59",     3614 => x"7A",     3615 => x"8E", 
    3616 => x"9A",     3617 => x"91",     3618 => x"7F",     3619 => x"6E",     3620 => x"5A",     3621 => x"5B",     3622 => x"6C",     3623 => x"82", 
    3624 => x"91",     3625 => x"83",     3626 => x"67",     3627 => x"3A",     3628 => x"1A",     3629 => x"1F",     3630 => x"3E",     3631 => x"80", 
    3632 => x"B9",     3633 => x"EA",     3634 => x"F0",     3635 => x"D0",     3636 => x"A3",     3637 => x"6A",     3638 => x"52",     3639 => x"4B", 
    3640 => x"66",     3641 => x"84",     3642 => x"95",     3643 => x"99",     3644 => x"7E",     3645 => x"62",     3646 => x"43",     3647 => x"3C", 
    3648 => x"4A",     3649 => x"60",     3650 => x"80",     3651 => x"90",     3652 => x"97",     3653 => x"8B",     3654 => x"7C",     3655 => x"6D", 
    3656 => x"5D",     3657 => x"60",     3658 => x"70",     3659 => x"84",     3660 => x"8E",     3661 => x"7F",     3662 => x"64",     3663 => x"39", 
    3664 => x"1C",     3665 => x"23",     3666 => x"41",     3667 => x"81",     3668 => x"B7",     3669 => x"E5",     3670 => x"E9",     3671 => x"CA", 
    3672 => x"9F",     3673 => x"6B",     3674 => x"58",     3675 => x"54",     3676 => x"6E",     3677 => x"87",     3678 => x"93",     3679 => x"92", 
    3680 => x"77",     3681 => x"5F",     3682 => x"45",     3683 => x"41",     3684 => x"4E",     3685 => x"63",     3686 => x"7F",     3687 => x"8C", 
    3688 => x"94",     3689 => x"89",     3690 => x"7C",     3691 => x"6F",     3692 => x"60",     3693 => x"5F",     3694 => x"6B",     3695 => x"7E", 
    3696 => x"8A",     3697 => x"80",     3698 => x"68",     3699 => x"41",     3700 => x"22",     3701 => x"26",     3702 => x"41",     3703 => x"7C", 
    3704 => x"B3",     3705 => x"DE",     3706 => x"E9",     3707 => x"CC",     3708 => x"A5",     3709 => x"72",     3710 => x"5A",     3711 => x"54", 
    3712 => x"68",     3713 => x"84",     3714 => x"91",     3715 => x"94",     3716 => x"7D",     3717 => x"64",     3718 => x"49",     3719 => x"3F", 
    3720 => x"49",     3721 => x"5B",     3722 => x"77",     3723 => x"88",     3724 => x"91",     3725 => x"8D",     3726 => x"81",     3727 => x"74", 
    3728 => x"63",     3729 => x"5B",     3730 => x"63",     3731 => x"75",     3732 => x"87",     3733 => x"85",     3734 => x"72",     3735 => x"52", 
    3736 => x"2D",     3737 => x"28",     3738 => x"3A",     3739 => x"6D",     3740 => x"A5",     3741 => x"D2",     3742 => x"E6",     3743 => x"CE", 
    3744 => x"A9",     3745 => x"78",     3746 => x"5B",     3747 => x"56",     3748 => x"65",     3749 => x"83",     3750 => x"90",     3751 => x"95", 
    3752 => x"81",     3753 => x"67",     3754 => x"4F",     3755 => x"41",     3756 => x"49",     3757 => x"58",     3758 => x"72",     3759 => x"85", 
    3760 => x"90",     3761 => x"92",     3762 => x"88",     3763 => x"7F",     3764 => x"6F",     3765 => x"62",     3766 => x"5A",     3767 => x"66", 
    3768 => x"78",     3769 => x"87",     3770 => x"86",     3771 => x"71",     3772 => x"53",     3773 => x"2F",     3774 => x"2F",     3775 => x"41", 
    3776 => x"74",     3777 => x"AA",     3778 => x"D1",     3779 => x"E0",     3780 => x"C3",     3781 => x"A1",     3782 => x"71",     3783 => x"5B", 
    3784 => x"59",     3785 => x"69",     3786 => x"84",     3787 => x"8E",     3788 => x"92",     3789 => x"7D",     3790 => x"66",     3791 => x"4F", 
    3792 => x"44",     3793 => x"4E",     3794 => x"5A",     3795 => x"73",     3796 => x"81",     3797 => x"8D",     3798 => x"8E",     3799 => x"85", 
    3800 => x"7D",     3801 => x"6B",     3802 => x"5E",     3803 => x"54",     3804 => x"62",     3805 => x"74",     3806 => x"87",     3807 => x"87", 
    3808 => x"72",     3809 => x"53",     3810 => x"2C",     3811 => x"2F",     3812 => x"40",     3813 => x"79",     3814 => x"AE",     3815 => x"D7", 
    3816 => x"E4",     3817 => x"C5",     3818 => x"A3",     3819 => x"71",     3820 => x"5E",     3821 => x"5D",     3822 => x"6F",     3823 => x"8C", 
    3824 => x"90",     3825 => x"92",     3826 => x"78",     3827 => x"61",     3828 => x"4C",     3829 => x"42",     3830 => x"4F",     3831 => x"59", 
    3832 => x"73",     3833 => x"80",     3834 => x"8C",     3835 => x"8C",     3836 => x"82",     3837 => x"7C",     3838 => x"6A",     3839 => x"60", 
    3840 => x"57",     3841 => x"66",     3842 => x"78",     3843 => x"89",     3844 => x"87",     3845 => x"70",     3846 => x"4F",     3847 => x"2A", 
    3848 => x"2F",     3849 => x"43",     3850 => x"7C",     3851 => x"B0",     3852 => x"D8",     3853 => x"E1",     3854 => x"C1",     3855 => x"9E", 
    3856 => x"6D",     3857 => x"5D",     3858 => x"5C",     3859 => x"71",     3860 => x"8A",     3861 => x"8E",     3862 => x"8D",     3863 => x"72", 
    3864 => x"5C",     3865 => x"48",     3866 => x"45",     3867 => x"52",     3868 => x"5E",     3869 => x"76",     3870 => x"80",     3871 => x"8B", 
    3872 => x"89",     3873 => x"83",     3874 => x"7E",     3875 => x"6E",     3876 => x"63",     3877 => x"5C",     3878 => x"6D",     3879 => x"7C", 
    3880 => x"8B",     3881 => x"81",     3882 => x"6A",     3883 => x"46",     3884 => x"28",     3885 => x"31",     3886 => x"49",     3887 => x"86", 
    3888 => x"B6",     3889 => x"DC",     3890 => x"DC",     3891 => x"BB",     3892 => x"96",     3893 => x"68",     3894 => x"5E",     3895 => x"5D", 
    3896 => x"75",     3897 => x"8A",     3898 => x"8F",     3899 => x"8D",     3900 => x"72",     3901 => x"60",     3902 => x"4A",     3903 => x"47", 
    3904 => x"51",     3905 => x"5E",     3906 => x"75",     3907 => x"80",     3908 => x"8C",     3909 => x"89",     3910 => x"84",     3911 => x"7A", 
    3912 => x"69",     3913 => x"5C",     3914 => x"5B",     3915 => x"6D",     3916 => x"7F",     3917 => x"8A",     3918 => x"7C",     3919 => x"63", 
    3920 => x"39",     3921 => x"29",     3922 => x"34",     3923 => x"5B",     3924 => x"99",     3925 => x"C5",     3926 => x"E5",     3927 => x"D3", 
    3928 => x"B2",     3929 => x"84",     3930 => x"61",     3931 => x"5E",     3932 => x"65",     3933 => x"83",     3934 => x"8F",     3935 => x"92", 
    3936 => x"82",     3937 => x"68",     3938 => x"54",     3939 => x"43",     3940 => x"4D",     3941 => x"58",     3942 => x"6B",     3943 => x"7D", 
    3944 => x"86",     3945 => x"8B",     3946 => x"84",     3947 => x"81",     3948 => x"74",     3949 => x"67",     3950 => x"5F",     3951 => x"67", 
    3952 => x"78",     3953 => x"88",     3954 => x"86",     3955 => x"71",     3956 => x"51",     3957 => x"2C",     3958 => x"2C",     3959 => x"40", 
    3960 => x"78",     3961 => x"AD",     3962 => x"D5",     3963 => x"E1",     3964 => x"C2",     3965 => x"A0",     3966 => x"6F",     3967 => x"5D", 
    3968 => x"5C",     3969 => x"6E",     3970 => x"87",     3971 => x"8C",     3972 => x"8C",     3973 => x"73",     3974 => x"5F",     3975 => x"4B", 
    3976 => x"44",     3977 => x"51",     3978 => x"5D",     3979 => x"75",     3980 => x"81",     3981 => x"8D",     3982 => x"8D",     3983 => x"86", 
    3984 => x"7F",     3985 => x"6F",     3986 => x"63",     3987 => x"5C",     3988 => x"6B",     3989 => x"7B",     3990 => x"89",     3991 => x"80", 
    3992 => x"69",     3993 => x"44",     3994 => x"27",     3995 => x"30",     3996 => x"4A",     3997 => x"86",     3998 => x"B6",     3999 => x"DC", 
    4000 => x"DB",     4001 => x"BB",     4002 => x"96",     4003 => x"69",     4004 => x"5E",     4005 => x"5F",     4006 => x"77",     4007 => x"8C", 
    4008 => x"90",     4009 => x"8B",     4010 => x"6E",     4011 => x"5C",     4012 => x"47",     4013 => x"48",     4014 => x"54",     4015 => x"63", 
    4016 => x"78",     4017 => x"82",     4018 => x"8C",     4019 => x"88",     4020 => x"84",     4021 => x"7A",     4022 => x"69",     4023 => x"5D", 
    4024 => x"5F",     4025 => x"6F",     4026 => x"80",     4027 => x"87",     4028 => x"76",     4029 => x"5A",     4030 => x"31",     4031 => x"27", 
    4032 => x"36",     4033 => x"64",     4034 => x"A0",     4035 => x"CB",     4036 => x"E5",     4037 => x"CF",     4038 => x"AE",     4039 => x"80", 
    4040 => x"62",     4041 => x"5E",     4042 => x"67",     4043 => x"82",     4044 => x"8C",     4045 => x"8F",     4046 => x"7F",     4047 => x"67", 
    4048 => x"54",     4049 => x"44",     4050 => x"4C",     4051 => x"55",     4052 => x"6A",     4053 => x"7B",     4054 => x"87",     4055 => x"8E", 
    4056 => x"86",     4057 => x"82",     4058 => x"72",     4059 => x"64",     4060 => x"5C",     4061 => x"68",     4062 => x"7A",     4063 => x"89", 
    4064 => x"85",     4065 => x"6F",     4066 => x"4A",     4067 => x"27",     4068 => x"2A",     4069 => x"44",     4070 => x"7F",     4071 => x"B4", 
    4072 => x"DB",     4073 => x"E0",     4074 => x"C0",     4075 => x"9A",     4076 => x"6C",     4077 => x"5D",     4078 => x"5C",     4079 => x"72", 
    4080 => x"8A",     4081 => x"8F",     4082 => x"8D",     4083 => x"73",     4084 => x"5D",     4085 => x"47",     4086 => x"42",     4087 => x"4E", 
    4088 => x"5D",     4089 => x"76",     4090 => x"85",     4091 => x"92",     4092 => x"91",     4093 => x"89",     4094 => x"7E",     4095 => x"6B", 
    4096 => x"5D",     4097 => x"5A",     4098 => x"6C",     4099 => x"7E",     4100 => x"8B",     4101 => x"7E",     4102 => x"65",     4103 => x"3B", 
    4104 => x"27",     4105 => x"30",     4106 => x"55",     4107 => x"94",     4108 => x"C2",     4109 => x"E4",     4110 => x"D7",     4111 => x"B5", 
    4112 => x"89",     4113 => x"63",     4114 => x"5C",     4115 => x"61",     4116 => x"7E",     4117 => x"8D",     4118 => x"92",     4119 => x"86", 
    4120 => x"6B",     4121 => x"57",     4122 => x"42",     4123 => x"47",     4124 => x"52",     4125 => x"66",     4126 => x"7D",     4127 => x"8A", 
    4128 => x"93",     4129 => x"8C",     4130 => x"84",     4131 => x"73",     4132 => x"62",     4133 => x"58",     4134 => x"60",     4135 => x"73", 
    4136 => x"85",     4137 => x"88",     4138 => x"76",     4139 => x"56",     4140 => x"2D",     4141 => x"27",     4142 => x"37",     4143 => x"6B", 
    4144 => x"A5",     4145 => x"D2",     4146 => x"E6",     4147 => x"CE",     4148 => x"AA",     4149 => x"7A",     4150 => x"61",     4151 => x"5D", 
    4152 => x"6C",     4153 => x"87",     4154 => x"90",     4155 => x"92",     4156 => x"7D",     4157 => x"65",     4158 => x"4D",     4159 => x"3F", 
    4160 => x"47",     4161 => x"52",     4162 => x"6C",     4163 => x"7F",     4164 => x"8E",     4165 => x"93",     4166 => x"8B",     4167 => x"81", 
    4168 => x"6D",     4169 => x"5C",     4170 => x"56",     4171 => x"66",     4172 => x"7A",     4173 => x"8A",     4174 => x"81",     4175 => x"69", 
    4176 => x"41",     4177 => x"25",     4178 => x"2A",     4179 => x"48",     4180 => x"84",     4181 => x"B8",     4182 => x"E1",     4183 => x"E4", 
    4184 => x"C7",     4185 => x"9E",     4186 => x"6E",     4187 => x"5C",     4188 => x"59",     4189 => x"72",     4190 => x"89",     4191 => x"92", 
    4192 => x"8F",     4193 => x"75",     4194 => x"5C",     4195 => x"41",     4196 => x"3D",     4197 => x"48",     4198 => x"5C",     4199 => x"78", 
    4200 => x"88",     4201 => x"93",     4202 => x"8F",     4203 => x"84",     4204 => x"75",     4205 => x"60",     4206 => x"5B",     4207 => x"66", 
    4208 => x"7A",     4209 => x"89",     4210 => x"80",     4211 => x"6A",     4212 => x"3F",     4213 => x"24",     4214 => x"27",     4215 => x"45", 
    4216 => x"81",     4217 => x"B7",     4218 => x"E3",     4219 => x"E7",     4220 => x"CD",     4221 => x"A2",     4222 => x"72",     4223 => x"5C", 
    4224 => x"58",     4225 => x"6E",     4226 => x"86",     4227 => x"92",     4228 => x"90",     4229 => x"78",     4230 => x"5E",     4231 => x"41", 
    4232 => x"39",     4233 => x"44",     4234 => x"58",     4235 => x"77",     4236 => x"8B",     4237 => x"98",     4238 => x"95",     4239 => x"87", 
    4240 => x"75",     4241 => x"5E",     4242 => x"59",     4243 => x"65",     4244 => x"79",     4245 => x"89",     4246 => x"7E",     4247 => x"68", 
    4248 => x"3D",     4249 => x"24",     4250 => x"28",     4251 => x"46",     4252 => x"82",     4253 => x"B7",     4254 => x"E3",     4255 => x"E6", 
    4256 => x"CE",     4257 => x"A6",     4258 => x"77",     4259 => x"61",     4260 => x"5B",     4261 => x"6F",     4262 => x"85",     4263 => x"8F", 
    4264 => x"8C",     4265 => x"74",     4266 => x"5C",     4267 => x"43",     4268 => x"3D",     4269 => x"48",     4270 => x"5B",     4271 => x"75", 
    4272 => x"87",     4273 => x"93",     4274 => x"92",     4275 => x"86",     4276 => x"76",     4277 => x"61",     4278 => x"60",     4279 => x"6B", 
    4280 => x"7A",     4281 => x"82",     4282 => x"73",     4283 => x"5D",     4284 => x"34",     4285 => x"25",     4286 => x"2D",     4287 => x"52", 
    4288 => x"8D",     4289 => x"BF",     4290 => x"E7",     4291 => x"E6",     4292 => x"CD",     4293 => x"A3",     4294 => x"77",     4295 => x"61", 
    4296 => x"5D",     4297 => x"70",     4298 => x"81",     4299 => x"87",     4300 => x"83",     4301 => x"6E",     4302 => x"5A",     4303 => x"47", 
    4304 => x"45",     4305 => x"4D",     4306 => x"5D",     4307 => x"75",     4308 => x"85",     4309 => x"92",     4310 => x"91",     4311 => x"86", 
    4312 => x"74",     4313 => x"62",     4314 => x"67",     4315 => x"6F",     4316 => x"7B",     4317 => x"75",     4318 => x"64",     4319 => x"46", 
    4320 => x"29",     4321 => x"2A",     4322 => x"3E",     4323 => x"6F",     4324 => x"A4",     4325 => x"D1",     4326 => x"E8",     4327 => x"DC", 
    4328 => x"BF",     4329 => x"95",     4330 => x"73",     4331 => x"64",     4332 => x"66",     4333 => x"76",     4334 => x"7D",     4335 => x"7F", 
    4336 => x"75",     4337 => x"61",     4338 => x"52",     4339 => x"47",     4340 => x"4A",     4341 => x"54",     4342 => x"66",     4343 => x"7D", 
    4344 => x"8B",     4345 => x"93",     4346 => x"8E",     4347 => x"80",     4348 => x"6D",     4349 => x"67",     4350 => x"6D",     4351 => x"75", 
    4352 => x"75",     4353 => x"68",     4354 => x"51",     4355 => x"33",     4356 => x"2A",     4357 => x"36",     4358 => x"59",     4359 => x"8C", 
    4360 => x"BC",     4361 => x"DD",     4362 => x"E2",     4363 => x"D0",     4364 => x"AF",     4365 => x"8B",     4366 => x"72",     4367 => x"68", 
    4368 => x"6C",     4369 => x"73",     4370 => x"74",     4371 => x"72",     4372 => x"67",     4373 => x"5B",     4374 => x"51",     4375 => x"4C", 
    4376 => x"51",     4377 => x"5B",     4378 => x"6D",     4379 => x"7E",     4380 => x"8A",     4381 => x"8E",     4382 => x"86",     4383 => x"77", 
    4384 => x"6F",     4385 => x"6F",     4386 => x"71",     4387 => x"6D",     4388 => x"62",     4389 => x"4F",     4390 => x"39",     4391 => x"34", 
    4392 => x"3E",     4393 => x"5C",     4394 => x"86",     4395 => x"AE",     4396 => x"CE",     4397 => x"D7",     4398 => x"CE",     4399 => x"B6", 
    4400 => x"99",     4401 => x"82",     4402 => x"73",     4403 => x"6E",     4404 => x"6D",     4405 => x"6C",     4406 => x"6B",     4407 => x"66", 
    4408 => x"5F",     4409 => x"58",     4410 => x"53",     4411 => x"53",     4412 => x"59",     4413 => x"68",     4414 => x"77",     4415 => x"82", 
    4416 => x"86",     4417 => x"81",     4418 => x"78",     4419 => x"76",     4420 => x"75",     4421 => x"74",     4422 => x"6D",     4423 => x"61", 
    4424 => x"50",     4425 => x"40",     4426 => x"40",     4427 => x"4B",     4428 => x"64",     4429 => x"85",     4430 => x"A4",     4431 => x"BC", 
    4432 => x"C6",     4433 => x"C4",     4434 => x"B7",     4435 => x"A3",     4436 => x"8F",     4437 => x"7F",     4438 => x"75",     4439 => x"6E", 
    4440 => x"6A",     4441 => x"68",     4442 => x"62",     4443 => x"5D",     4444 => x"57",     4445 => x"53",     4446 => x"53",     4447 => x"59", 
    4448 => x"64",     4449 => x"70",     4450 => x"7A",     4451 => x"7E",     4452 => x"7C",     4453 => x"7C",     4454 => x"7A",     4455 => x"77", 
    4456 => x"70",     4457 => x"64",     4458 => x"57",     4459 => x"4B",     4460 => x"4A",     4461 => x"51",     4462 => x"62",     4463 => x"7A", 
    4464 => x"91",     4465 => x"A5",     4466 => x"B1",     4467 => x"B5",     4468 => x"B2",     4469 => x"A8",     4470 => x"9C",     4471 => x"91", 
    4472 => x"88",     4473 => x"80",     4474 => x"77",     4475 => x"70",     4476 => x"67",     4477 => x"5D",     4478 => x"57",     4479 => x"53", 
    4480 => x"52",     4481 => x"56",     4482 => x"5C",     4483 => x"64",     4484 => x"6C",     4485 => x"70",     4486 => x"75",     4487 => x"7B", 
    4488 => x"7E",     4489 => x"7C",     4490 => x"74",     4491 => x"68",     4492 => x"5A",     4493 => x"53",     4494 => x"56",     4495 => x"60", 
    4496 => x"70",     4497 => x"81",     4498 => x"91",     4499 => x"9B",     4500 => x"A2",     4501 => x"A3",     4502 => x"A1",     4503 => x"9E", 
    4504 => x"9C",     4505 => x"98",     4506 => x"92",     4507 => x"89",     4508 => x"7E",     4509 => x"73",     4510 => x"68",     4511 => x"5F", 
    4512 => x"5A",     4513 => x"57",     4514 => x"55",     4515 => x"56",     4516 => x"59",     4517 => x"5C",     4518 => x"5E",     4519 => x"67", 
    4520 => x"6F",     4521 => x"74",     4522 => x"75",     4523 => x"72",     4524 => x"6A",     4525 => x"63",     4526 => x"61",     4527 => x"64", 
    4528 => x"6A",     4529 => x"74",     4530 => x"7F",     4531 => x"88",     4532 => x"90",     4533 => x"95",     4534 => x"9A",     4535 => x"9E", 
    4536 => x"A0",     4537 => x"A0",     4538 => x"9B",     4539 => x"93",     4540 => x"8A",     4541 => x"81",     4542 => x"79",     4543 => x"71", 
    4544 => x"6A",     4545 => x"63",     4546 => x"5D",     4547 => x"59",     4548 => x"56",     4549 => x"55",     4550 => x"55",     4551 => x"5A", 
    4552 => x"60",     4553 => x"63",     4554 => x"66",     4555 => x"66",     4556 => x"64",     4557 => x"64",     4558 => x"68",     4559 => x"6E", 
    4560 => x"75",     4561 => x"7C",     4562 => x"81",     4563 => x"84",     4564 => x"88",     4565 => x"8E",     4566 => x"96",     4567 => x"9D", 
    4568 => x"A2",     4569 => x"A3",     4570 => x"9E",     4571 => x"97",     4572 => x"8F",     4573 => x"87",     4574 => x"7F",     4575 => x"76", 
    4576 => x"6E",     4577 => x"65",     4578 => x"5D",     4579 => x"57",     4580 => x"55",     4581 => x"53",     4582 => x"53",     4583 => x"56", 
    4584 => x"57",     4585 => x"59",     4586 => x"5B",     4587 => x"5F",     4588 => x"62",     4589 => x"67",     4590 => x"6D",     4591 => x"73", 
    4592 => x"79",     4593 => x"7F",     4594 => x"85",     4595 => x"8A",     4596 => x"90",     4597 => x"96",     4598 => x"9C",     4599 => x"A1", 
    4600 => x"A3",     4601 => x"A2",     4602 => x"9F",     4603 => x"99",     4604 => x"91",     4605 => x"87",     4606 => x"7D",     4607 => x"71", 
    4608 => x"66",     4609 => x"5C",     4610 => x"53",     4611 => x"4F",     4612 => x"4D",     4613 => x"4D",     4614 => x"4F",     4615 => x"53", 
    4616 => x"56",     4617 => x"59",     4618 => x"5D",     4619 => x"63",     4620 => x"68",     4621 => x"6E",     4622 => x"73",     4623 => x"7A", 
    4624 => x"80",     4625 => x"88",     4626 => x"90",     4627 => x"96",     4628 => x"9C",     4629 => x"A1",     4630 => x"A4",     4631 => x"A4", 
    4632 => x"A2",     4633 => x"9D",     4634 => x"96",     4635 => x"8C",     4636 => x"82",     4637 => x"76",     4638 => x"69",     4639 => x"5E", 
    4640 => x"55",     4641 => x"4D",     4642 => x"48",     4643 => x"48",     4644 => x"4A",     4645 => x"4E",     4646 => x"53",     4647 => x"58", 
    4648 => x"5E",     4649 => x"64",     4650 => x"69",     4651 => x"70",     4652 => x"77",     4653 => x"7E",     4654 => x"85",     4655 => x"8C", 
    4656 => x"92",     4657 => x"98",     4658 => x"9D",     4659 => x"A1",     4660 => x"A4",     4661 => x"A4",     4662 => x"A2",     4663 => x"9C", 
    4664 => x"94",     4665 => x"8A",     4666 => x"7D",     4667 => x"71",     4668 => x"64",     4669 => x"5A",     4670 => x"52",     4671 => x"4C", 
    4672 => x"48",     4673 => x"47",     4674 => x"4A",     4675 => x"4E",     4676 => x"54",     4677 => x"5A",     4678 => x"61",     4679 => x"67", 
    4680 => x"6E",     4681 => x"75",     4682 => x"7C",     4683 => x"82",     4684 => x"88",     4685 => x"8E",     4686 => x"94",     4687 => x"99", 
    4688 => x"9D",     4689 => x"A0",     4690 => x"A1",     4691 => x"A0",     4692 => x"9B",     4693 => x"95",     4694 => x"8C",     4695 => x"83", 
    4696 => x"78",     4697 => x"6D",     4698 => x"62",     4699 => x"59",     4700 => x"52",     4701 => x"4E",     4702 => x"4B",     4703 => x"4B", 
    4704 => x"4C",     4705 => x"50",     4706 => x"55",     4707 => x"5B",     4708 => x"62",     4709 => x"69",     4710 => x"70",     4711 => x"77", 
    4712 => x"7E",     4713 => x"86",     4714 => x"8D",     4715 => x"93",     4716 => x"98",     4717 => x"9C",     4718 => x"9E",     4719 => x"9E", 
    4720 => x"9E",     4721 => x"9B",     4722 => x"96",     4723 => x"90",     4724 => x"89",     4725 => x"80",     4726 => x"77",     4727 => x"6D", 
    4728 => x"64",     4729 => x"5C",     4730 => x"55",     4731 => x"51",     4732 => x"4F",     4733 => x"4E",     4734 => x"50",     4735 => x"52", 
    4736 => x"56",     4737 => x"5A",     4738 => x"61",     4739 => x"68",     4740 => x"6F",     4741 => x"75",     4742 => x"7B",     4743 => x"81", 
    4744 => x"88",     4745 => x"8F",     4746 => x"95",     4747 => x"9A",     4748 => x"9C",     4749 => x"9D",     4750 => x"9C",     4751 => x"9A", 
    4752 => x"96",     4753 => x"90",     4754 => x"89",     4755 => x"80",     4756 => x"77",     4757 => x"6F",     4758 => x"66",     4759 => x"60", 
    4760 => x"5A",     4761 => x"55",     4762 => x"52",     4763 => x"51",     4764 => x"52",     4765 => x"54",     4766 => x"56",     4767 => x"5A", 
    4768 => x"5F",     4769 => x"64",     4770 => x"6B",     4771 => x"71",     4772 => x"78",     4773 => x"7E",     4774 => x"85",     4775 => x"8B", 
    4776 => x"90",     4777 => x"94",     4778 => x"98",     4779 => x"99",     4780 => x"9A",     4781 => x"99",     4782 => x"97",     4783 => x"93", 
    4784 => x"8E",     4785 => x"88",     4786 => x"80",     4787 => x"77",     4788 => x"6F",     4789 => x"66",     4790 => x"60",     4791 => x"5C", 
    4792 => x"59",     4793 => x"58",     4794 => x"57",     4795 => x"56",     4796 => x"57",     4797 => x"59",     4798 => x"5D",     4799 => x"61", 
    4800 => x"67",     4801 => x"6D",     4802 => x"73",     4803 => x"79",     4804 => x"7E",     4805 => x"82",     4806 => x"86",     4807 => x"8B", 
    4808 => x"8F",     4809 => x"92",     4810 => x"94",     4811 => x"94",     4812 => x"93",     4813 => x"92",     4814 => x"8F",     4815 => x"8B", 
    4816 => x"87",     4817 => x"80",     4818 => x"7A",     4819 => x"73",     4820 => x"6D",     4821 => x"67",     4822 => x"61",     4823 => x"5D", 
    4824 => x"5A",     4825 => x"58",     4826 => x"57",     4827 => x"57",     4828 => x"59",     4829 => x"5D",     4830 => x"60",     4831 => x"64", 
    4832 => x"69",     4833 => x"6F",     4834 => x"75",     4835 => x"7A",     4836 => x"81",     4837 => x"86",     4838 => x"8A",     4839 => x"8E", 
    4840 => x"90",     4841 => x"92",     4842 => x"91",     4843 => x"90",     4844 => x"8F",     4845 => x"8D",     4846 => x"8B",     4847 => x"88", 
    4848 => x"83",     4849 => x"7F",     4850 => x"79",     4851 => x"73",     4852 => x"6E",     4853 => x"6A",     4854 => x"67",     4855 => x"64", 
    4856 => x"62",     4857 => x"61",     4858 => x"5F",     4859 => x"5D",     4860 => x"5D",     4861 => x"5E",     4862 => x"61",     4863 => x"66", 
    4864 => x"6B",     4865 => x"6F",     4866 => x"73",     4867 => x"78",     4868 => x"7A",     4869 => x"7F",     4870 => x"83",     4871 => x"89", 
    4872 => x"8B",     4873 => x"8E",     4874 => x"8F",     4875 => x"90",     4876 => x"8F",     4877 => x"8C",     4878 => x"89",     4879 => x"85", 
    4880 => x"80",     4881 => x"7C",     4882 => x"78",     4883 => x"74",     4884 => x"70",     4885 => x"6B",     4886 => x"66",     4887 => x"62", 
    4888 => x"60",     4889 => x"5F",     4890 => x"5F",     4891 => x"60",     4892 => x"62",     4893 => x"63",     4894 => x"65",     4895 => x"66", 
    4896 => x"6A",     4897 => x"6D",     4898 => x"72",     4899 => x"77",     4900 => x"7B",     4901 => x"7E",     4902 => x"82",     4903 => x"87", 
    4904 => x"88",     4905 => x"8B",     4906 => x"8C",     4907 => x"8D",     4908 => x"8C",     4909 => x"8B",     4910 => x"8A",     4911 => x"88", 
    4912 => x"85",     4913 => x"81",     4914 => x"7C",     4915 => x"77",     4916 => x"72",     4917 => x"6E",     4918 => x"6B",     4919 => x"67", 
    4920 => x"64",     4921 => x"62",     4922 => x"60",     4923 => x"5F",     4924 => x"61",     4925 => x"63",     4926 => x"64",     4927 => x"67", 
    4928 => x"6A",     4929 => x"6D",     4930 => x"70",     4931 => x"74",     4932 => x"77",     4933 => x"7A",     4934 => x"7E",     4935 => x"81", 
    4936 => x"84",     4937 => x"87",     4938 => x"8A",     4939 => x"8B",     4940 => x"8A",     4941 => x"89",     4942 => x"87",     4943 => x"86", 
    4944 => x"83",     4945 => x"81",     4946 => x"7D",     4947 => x"79",     4948 => x"75",     4949 => x"71",     4950 => x"6C",     4951 => x"68", 
    4952 => x"67",     4953 => x"65",     4954 => x"65",     4955 => x"65",     4956 => x"66",     4957 => x"66",     4958 => x"68",     4959 => x"69", 
    4960 => x"6B",     4961 => x"6D",     4962 => x"6E",     4963 => x"71",     4964 => x"73",     4965 => x"76",     4966 => x"7A",     4967 => x"7C", 
    4968 => x"81",     4969 => x"84",     4970 => x"86",     4971 => x"87",     4972 => x"88",     4973 => x"89",     4974 => x"89",     4975 => x"88", 
    4976 => x"85",     4977 => x"82",     4978 => x"7E",     4979 => x"7A",     4980 => x"75",     4981 => x"73",     4982 => x"70",     4983 => x"6D", 
    4984 => x"6B",     4985 => x"6A",     4986 => x"67",     4987 => x"67",     4988 => x"68",     4989 => x"69",     4990 => x"6A",     4991 => x"6A", 
    4992 => x"6C",     4993 => x"6C",     4994 => x"6C",     4995 => x"6D",     4996 => x"6F",     4997 => x"71",     4998 => x"73",     4999 => x"77", 
    5000 => x"79",     5001 => x"7F",     5002 => x"83",     5003 => x"87",     5004 => x"88",     5005 => x"89",     5006 => x"88",     5007 => x"88", 
    5008 => x"87",     5009 => x"86",     5010 => x"83",     5011 => x"7F",     5012 => x"7A",     5013 => x"76",     5014 => x"73",     5015 => x"70", 
    5016 => x"6F",     5017 => x"6C",     5018 => x"6B",     5019 => x"6A",     5020 => x"6A",     5021 => x"6B",     5022 => x"6C",     5023 => x"6C", 
    5024 => x"6D",     5025 => x"6D",     5026 => x"6E",     5027 => x"6E",     5028 => x"6E",     5029 => x"6F",     5030 => x"71",     5031 => x"72", 
    5032 => x"74",     5033 => x"77",     5034 => x"7B",     5035 => x"7E",     5036 => x"81",     5037 => x"84",     5038 => x"85",     5039 => x"87", 
    5040 => x"88",     5041 => x"86",     5042 => x"86",     5043 => x"83",     5044 => x"80",     5045 => x"7C",     5046 => x"79",     5047 => x"76", 
    5048 => x"72",     5049 => x"6F",     5050 => x"6D",     5051 => x"6B",     5052 => x"67",     5053 => x"66",     5054 => x"67",     5055 => x"68", 
    5056 => x"6B",     5057 => x"6B",     5058 => x"6C",     5059 => x"6B",     5060 => x"6C",     5061 => x"6E",     5062 => x"71",     5063 => x"74", 
    5064 => x"76",     5065 => x"77",     5066 => x"79",     5067 => x"7D",     5068 => x"80",     5069 => x"83",     5070 => x"83",     5071 => x"84", 
    5072 => x"85",     5073 => x"86",     5074 => x"86",     5075 => x"85",     5076 => x"84",     5077 => x"7F",     5078 => x"7B",     5079 => x"76", 
    5080 => x"73",     5081 => x"71",     5082 => x"71",     5083 => x"70",     5084 => x"6F",     5085 => x"6B",     5086 => x"6A",     5087 => x"6A", 
    5088 => x"6B",     5089 => x"6B",     5090 => x"68",     5091 => x"67",     5092 => x"67",     5093 => x"6B",     5094 => x"6E",     5095 => x"72", 
    5096 => x"73",     5097 => x"76",     5098 => x"7C",     5099 => x"7F",     5100 => x"83",     5101 => x"82",     5102 => x"83",     5103 => x"81", 
    5104 => x"84",     5105 => x"84",     5106 => x"85",     5107 => x"82",     5108 => x"81",     5109 => x"80",     5110 => x"7D",     5111 => x"79", 
    5112 => x"73",     5113 => x"6F",     5114 => x"6E",     5115 => x"70",     5116 => x"6E",     5117 => x"6D",     5118 => x"69",     5119 => x"6B", 
    5120 => x"6D",     5121 => x"71",     5122 => x"70",     5123 => x"70",     5124 => x"6D",     5125 => x"6C",     5126 => x"6E",     5127 => x"70", 
    5128 => x"74",     5129 => x"76",     5130 => x"7A",     5131 => x"7C",     5132 => x"7F",     5133 => x"80",     5134 => x"83",     5135 => x"84", 
    5136 => x"87",     5137 => x"87",     5138 => x"84",     5139 => x"81",     5140 => x"7F",     5141 => x"7F",     5142 => x"7D",     5143 => x"79", 
    5144 => x"72",     5145 => x"6E",     5146 => x"6C",     5147 => x"6E",     5148 => x"70",     5149 => x"6E",     5150 => x"6C",     5151 => x"68", 
    5152 => x"69",     5153 => x"6B",     5154 => x"6F",     5155 => x"6D",     5156 => x"6C",     5157 => x"6A",     5158 => x"6B",     5159 => x"6D", 
    5160 => x"70",     5161 => x"75",     5162 => x"78",     5163 => x"7C",     5164 => x"7F",     5165 => x"83",     5166 => x"84",     5167 => x"85", 
    5168 => x"85",     5169 => x"86",     5170 => x"87",     5171 => x"87",     5172 => x"86",     5173 => x"80",     5174 => x"7D",     5175 => x"75", 
    5176 => x"72",     5177 => x"70",     5178 => x"6F",     5179 => x"70",     5180 => x"6E",     5181 => x"6B",     5182 => x"69",     5183 => x"6A", 
    5184 => x"6D",     5185 => x"71",     5186 => x"71",     5187 => x"6F",     5188 => x"6B",     5189 => x"6A",     5190 => x"6A",     5191 => x"6D", 
    5192 => x"70",     5193 => x"71",     5194 => x"76",     5195 => x"77",     5196 => x"7D",     5197 => x"80",     5198 => x"84",     5199 => x"86", 
    5200 => x"88",     5201 => x"88",     5202 => x"89",     5203 => x"88",     5204 => x"84",     5205 => x"81",     5206 => x"7B",     5207 => x"7A", 
    5208 => x"77",     5209 => x"75",     5210 => x"70",     5211 => x"6D",     5212 => x"6A",     5213 => x"69",     5214 => x"6C",     5215 => x"6F", 
    5216 => x"6D",     5217 => x"6A",     5218 => x"67",     5219 => x"66",     5220 => x"69",     5221 => x"6D",     5222 => x"70",     5223 => x"71", 
    5224 => x"70",     5225 => x"72",     5226 => x"76",     5227 => x"7B",     5228 => x"82",     5229 => x"86",     5230 => x"87",     5231 => x"87", 
    5232 => x"86",     5233 => x"87",     5234 => x"87",     5235 => x"86",     5236 => x"84",     5237 => x"80",     5238 => x"7D",     5239 => x"7A", 
    5240 => x"77",     5241 => x"74",     5242 => x"71",     5243 => x"6F",     5244 => x"6F",     5245 => x"6F",     5246 => x"6E",     5247 => x"6A", 
    5248 => x"6B",     5249 => x"6B",     5250 => x"6C",     5251 => x"69",     5252 => x"68",     5253 => x"66",     5254 => x"67",     5255 => x"6C", 
    5256 => x"71",     5257 => x"77",     5258 => x"78",     5259 => x"7D",     5260 => x"80",     5261 => x"87",     5262 => x"88",     5263 => x"8A", 
    5264 => x"88",     5265 => x"88",     5266 => x"88",     5267 => x"88",     5268 => x"84",     5269 => x"7C",     5270 => x"77",     5271 => x"71", 
    5272 => x"71",     5273 => x"6E",     5274 => x"6E",     5275 => x"69",     5276 => x"68",     5277 => x"66",     5278 => x"6A",     5279 => x"6A", 
    5280 => x"6B",     5281 => x"6A",     5282 => x"68",     5283 => x"6C",     5284 => x"6C",     5285 => x"6E",     5286 => x"6A",     5287 => x"6C", 
    5288 => x"6C",     5289 => x"71",     5290 => x"79",     5291 => x"7F",     5292 => x"85",     5293 => x"85",     5294 => x"88",     5295 => x"89", 
    5296 => x"8A",     5297 => x"88",     5298 => x"83",     5299 => x"7F",     5300 => x"7E",     5301 => x"7D",     5302 => x"7A",     5303 => x"76", 
    5304 => x"71",     5305 => x"6C",     5306 => x"6C",     5307 => x"6B",     5308 => x"6B",     5309 => x"6B",     5310 => x"6A",     5311 => x"6C", 
    5312 => x"69",     5313 => x"67",     5314 => x"67",     5315 => x"67",     5316 => x"69",     5317 => x"6F",     5318 => x"70",     5319 => x"73", 
    5320 => x"75",     5321 => x"77",     5322 => x"7D",     5323 => x"82",     5324 => x"87",     5325 => x"89",     5326 => x"88",     5327 => x"86", 
    5328 => x"86",     5329 => x"86",     5330 => x"87",     5331 => x"82",     5332 => x"7E",     5333 => x"79",     5334 => x"77",     5335 => x"75", 
    5336 => x"73",     5337 => x"71",     5338 => x"6E",     5339 => x"71",     5340 => x"6F",     5341 => x"71",     5342 => x"70",     5343 => x"6E", 
    5344 => x"6C",     5345 => x"6E",     5346 => x"71",     5347 => x"72",     5348 => x"74",     5349 => x"73",     5350 => x"78",     5351 => x"7B", 
    5352 => x"82",     5353 => x"87",     5354 => x"8A",     5355 => x"88",     5356 => x"88",     5357 => x"87",     5358 => x"88",     5359 => x"89", 
    5360 => x"86",     5361 => x"83",     5362 => x"7B",     5363 => x"77",     5364 => x"71",     5365 => x"71",     5366 => x"6C",     5367 => x"6B", 
    5368 => x"67",     5369 => x"64",     5370 => x"62",     5371 => x"61",     5372 => x"65",     5373 => x"64",     5374 => x"67",     5375 => x"60", 
    5376 => x"5F",     5377 => x"5B",     5378 => x"5E",     5379 => x"60",     5380 => x"61",     5381 => x"67",     5382 => x"66",     5383 => x"71", 
    5384 => x"73",     5385 => x"7E",     5386 => x"80",     5387 => x"84",     5388 => x"83",     5389 => x"80",     5390 => x"81",     5391 => x"7F", 
    5392 => x"7F",     5393 => x"7A",     5394 => x"77",     5395 => x"70",     5396 => x"6F",     5397 => x"6C",     5398 => x"6C",     5399 => x"69", 
    5400 => x"68",     5401 => x"6B",     5402 => x"6B",     5403 => x"72",     5404 => x"6F",     5405 => x"6E",     5406 => x"66",     5407 => x"6B", 
    5408 => x"6C",     5409 => x"72",     5410 => x"75",     5411 => x"76",     5412 => x"7A",     5413 => x"7A",     5414 => x"82",     5415 => x"86", 
    5416 => x"8E",     5417 => x"8A",     5418 => x"8D",     5419 => x"8D",     5420 => x"92",     5421 => x"91",     5422 => x"90",     5423 => x"8B", 
    5424 => x"88",     5425 => x"88",     5426 => x"84",     5427 => x"81",     5428 => x"7A",     5429 => x"78",     5430 => x"75",     5431 => x"78", 
    5432 => x"7A",     5433 => x"7B",     5434 => x"79",     5435 => x"73",     5436 => x"75",     5437 => x"72",     5438 => x"75",     5439 => x"74", 
    5440 => x"75",     5441 => x"77",     5442 => x"78",     5443 => x"7B",     5444 => x"7B",     5445 => x"83",     5446 => x"87",     5447 => x"8C", 
    5448 => x"8C",     5449 => x"8E",     5450 => x"8F",     5451 => x"8E",     5452 => x"8E",     5453 => x"88",     5454 => x"88",     5455 => x"82", 
    5456 => x"80",     5457 => x"7B",     5458 => x"77",     5459 => x"72",     5460 => x"6F",     5461 => x"70",     5462 => x"70",     5463 => x"6D", 
    5464 => x"6B",     5465 => x"68",     5466 => x"6B",     5467 => x"6D",     5468 => x"6C",     5469 => x"67",     5470 => x"62",     5471 => x"65", 
    5472 => x"6A",     5473 => x"6D",     5474 => x"71",     5475 => x"6F",     5476 => x"72",     5477 => x"77",     5478 => x"7E",     5479 => x"82", 
    5480 => x"80",     5481 => x"7D",     5482 => x"7C",     5483 => x"80",     5484 => x"7F",     5485 => x"7D",     5486 => x"74",     5487 => x"6E", 
    5488 => x"69",     5489 => x"69",     5490 => x"69",     5491 => x"68",     5492 => x"67",     5493 => x"61",     5494 => x"63",     5495 => x"63", 
    5496 => x"6A",     5497 => x"69",     5498 => x"67",     5499 => x"64",     5500 => x"64",     5501 => x"64",     5502 => x"67",     5503 => x"66", 
    5504 => x"66",     5505 => x"6A",     5506 => x"6F",     5507 => x"75",     5508 => x"78",     5509 => x"7A",     5510 => x"7B",     5511 => x"7E", 
    5512 => x"7F",     5513 => x"80",     5514 => x"7D",     5515 => x"77",     5516 => x"75",     5517 => x"74",     5518 => x"74",     5519 => x"71", 
    5520 => x"6E",     5521 => x"6D",     5522 => x"6C",     5523 => x"6A",     5524 => x"6A",     5525 => x"6B",     5526 => x"6A",     5527 => x"6C", 
    5528 => x"6B",     5529 => x"6A",     5530 => x"69",     5531 => x"67",     5532 => x"6B",     5533 => x"6E",     5534 => x"74",     5535 => x"75", 
    5536 => x"78",     5537 => x"77",     5538 => x"7D",     5539 => x"81",     5540 => x"85",     5541 => x"86",     5542 => x"86",     5543 => x"86", 
    5544 => x"85",     5545 => x"83",     5546 => x"81",     5547 => x"7D",     5548 => x"7A",     5549 => x"7A",     5550 => x"77",     5551 => x"76", 
    5552 => x"72",     5553 => x"74",     5554 => x"74",     5555 => x"75",     5556 => x"78",     5557 => x"75",     5558 => x"74",     5559 => x"73", 
    5560 => x"74",     5561 => x"72",     5562 => x"72",     5563 => x"6E",     5564 => x"70",     5565 => x"72",     5566 => x"78",     5567 => x"7A", 
    5568 => x"7E",     5569 => x"80",     5570 => x"83",     5571 => x"86",     5572 => x"89",     5573 => x"8B",     5574 => x"88",     5575 => x"88", 
    5576 => x"82",     5577 => x"82",     5578 => x"7E",     5579 => x"7C",     5580 => x"7B",     5581 => x"79",     5582 => x"79",     5583 => x"77", 
    5584 => x"75",     5585 => x"73",     5586 => x"75",     5587 => x"71",     5588 => x"77",     5589 => x"72",     5590 => x"71",     5591 => x"6F", 
    5592 => x"6F",     5593 => x"71",     5594 => x"72",     5595 => x"74",     5596 => x"73",     5597 => x"74",     5598 => x"78",     5599 => x"7A", 
    5600 => x"7D",     5601 => x"7F",     5602 => x"80",     5603 => x"81",     5604 => x"83",     5605 => x"84",     5606 => x"84",     5607 => x"83", 
    5608 => x"7F",     5609 => x"7B",     5610 => x"78",     5611 => x"76",     5612 => x"77",     5613 => x"75",     5614 => x"73",     5615 => x"6F", 
    5616 => x"70",     5617 => x"71",     5618 => x"73",     5619 => x"72",     5620 => x"74",     5621 => x"6F",     5622 => x"6F",     5623 => x"72", 
    5624 => x"73",     5625 => x"73",     5626 => x"71",     5627 => x"71",     5628 => x"73",     5629 => x"77",     5630 => x"7A",     5631 => x"7D", 
    5632 => x"7F",     5633 => x"81",     5634 => x"80",     5635 => x"7E",     5636 => x"7C",     5637 => x"79",     5638 => x"79",     5639 => x"78", 
    5640 => x"78",     5641 => x"75",     5642 => x"71",     5643 => x"70",     5644 => x"71",     5645 => x"75",     5646 => x"72",     5647 => x"72", 
    5648 => x"6F",     5649 => x"70",     5650 => x"70",     5651 => x"72",     5652 => x"6F",     5653 => x"6D",     5654 => x"6F",     5655 => x"6F", 
    5656 => x"72",     5657 => x"74",     5658 => x"76",     5659 => x"76",     5660 => x"78",     5661 => x"7C",     5662 => x"7F",     5663 => x"81", 
    5664 => x"80",     5665 => x"7F",     5666 => x"7E",     5667 => x"7D",     5668 => x"7B",     5669 => x"77",     5670 => x"77",     5671 => x"76", 
    5672 => x"78",     5673 => x"75",     5674 => x"71",     5675 => x"71",     5676 => x"6F",     5677 => x"74",     5678 => x"72",     5679 => x"74", 
    5680 => x"6F",     5681 => x"71",     5682 => x"6E",     5683 => x"6D",     5684 => x"6C",     5685 => x"6A",     5686 => x"6C",     5687 => x"6B", 
    5688 => x"73",     5689 => x"6E",     5690 => x"73",     5691 => x"70",     5692 => x"74",     5693 => x"77",     5694 => x"7A",     5695 => x"78", 
    5696 => x"75",     5697 => x"75",     5698 => x"73",     5699 => x"77",     5700 => x"74",     5701 => x"76",     5702 => x"71",     5703 => x"72", 
    5704 => x"72",     5705 => x"75",     5706 => x"75",     5707 => x"72",     5708 => x"71",     5709 => x"71",     5710 => x"74",     5711 => x"73", 
    5712 => x"73",     5713 => x"6E",     5714 => x"6F",     5715 => x"70",     5716 => x"75",     5717 => x"75",     5718 => x"74",     5719 => x"73", 
    5720 => x"74",     5721 => x"7A",     5722 => x"79",     5723 => x"7C",     5724 => x"79",     5725 => x"7E",     5726 => x"7E",     5727 => x"7E", 
    5728 => x"7B",     5729 => x"76",     5730 => x"7A",     5731 => x"78",     5732 => x"7B",     5733 => x"77",     5734 => x"76",     5735 => x"72", 
    5736 => x"75",     5737 => x"77",     5738 => x"77",     5739 => x"77",     5740 => x"74",     5741 => x"78",     5742 => x"78",     5743 => x"7A", 
    5744 => x"75",     5745 => x"73",     5746 => x"72",     5747 => x"75",     5748 => x"77",     5749 => x"77",     5750 => x"76",     5751 => x"78", 
    5752 => x"7A",     5753 => x"7D",     5754 => x"7F",     5755 => x"7E",     5756 => x"7D",     5757 => x"80",     5758 => x"80",     5759 => x"81", 
    5760 => x"7F",     5761 => x"7B",     5762 => x"7D",     5763 => x"7C",     5764 => x"7D",     5765 => x"78",     5766 => x"79",     5767 => x"77", 
    5768 => x"7B",     5769 => x"7C",     5770 => x"7A",     5771 => x"7C",     5772 => x"7A",     5773 => x"7C",     5774 => x"77",     5775 => x"7B", 
    5776 => x"75",     5777 => x"76",     5778 => x"78",     5779 => x"78",     5780 => x"7A",     5781 => x"78",     5782 => x"75",     5783 => x"76", 
    5784 => x"79",     5785 => x"7A",     5786 => x"7D",     5787 => x"7E",     5788 => x"7E",     5789 => x"7D",     5790 => x"7E",     5791 => x"7B", 
    5792 => x"7C",     5793 => x"7A",     5794 => x"77",     5795 => x"77",     5796 => x"76",     5797 => x"77",     5798 => x"75",     5799 => x"78", 
    5800 => x"76",     5801 => x"79",     5802 => x"75",     5803 => x"77",     5804 => x"74",     5805 => x"73",     5806 => x"71",     5807 => x"71", 
    5808 => x"70",     5809 => x"73",     5810 => x"75",     5811 => x"72",     5812 => x"72",     5813 => x"6E",     5814 => x"70",     5815 => x"71", 
    5816 => x"75",     5817 => x"75",     5818 => x"73",     5819 => x"75",     5820 => x"73",     5821 => x"77",     5822 => x"74",     5823 => x"73", 
    5824 => x"72",     5825 => x"78",     5826 => x"78",     5827 => x"76",     5828 => x"73",     5829 => x"71",     5830 => x"71",     5831 => x"72", 
    5832 => x"76",     5833 => x"6E",     5834 => x"6E",     5835 => x"69",     5836 => x"6E",     5837 => x"6F",     5838 => x"70",     5839 => x"6B", 
    5840 => x"6B",     5841 => x"6D",     5842 => x"6E",     5843 => x"73",     5844 => x"6D",     5845 => x"70",     5846 => x"6D",     5847 => x"74", 
    5848 => x"74",     5849 => x"7A",     5850 => x"76",     5851 => x"73",     5852 => x"74",     5853 => x"74",     5854 => x"7A",     5855 => x"76", 
    5856 => x"77",     5857 => x"73",     5858 => x"77",     5859 => x"78",     5860 => x"7A",     5861 => x"78",     5862 => x"75",     5863 => x"77", 
    5864 => x"74",     5865 => x"77",     5866 => x"75",     5867 => x"73",     5868 => x"71",     5869 => x"6F",     5870 => x"72",     5871 => x"73", 
    5872 => x"74",     5873 => x"72",     5874 => x"72",     5875 => x"74",     5876 => x"77",     5877 => x"77",     5878 => x"77",     5879 => x"78", 
    5880 => x"76",     5881 => x"7D",     5882 => x"7D",     5883 => x"7E",     5884 => x"7B",     5885 => x"7A",     5886 => x"7A",     5887 => x"7B", 
    5888 => x"7B",     5889 => x"7A",     5890 => x"78",     5891 => x"7A",     5892 => x"7B",     5893 => x"7A",     5894 => x"7C",     5895 => x"76", 
    5896 => x"78",     5897 => x"77",     5898 => x"77",     5899 => x"77",     5900 => x"75",     5901 => x"74",     5902 => x"75",     5903 => x"77", 
    5904 => x"75",     5905 => x"75",     5906 => x"72",     5907 => x"72",     5908 => x"74",     5909 => x"77",     5910 => x"78",     5911 => x"76", 
    5912 => x"77",     5913 => x"78",     5914 => x"7B",     5915 => x"7E",     5916 => x"7A",     5917 => x"77",     5918 => x"78",     5919 => x"7A", 
    5920 => x"7A",     5921 => x"7A",     5922 => x"75",     5923 => x"76",     5924 => x"77",     5925 => x"7A",     5926 => x"78",     5927 => x"75", 
    5928 => x"73",     5929 => x"75",     5930 => x"75",     5931 => x"77",     5932 => x"74",     5933 => x"72",     5934 => x"74",     5935 => x"75", 
    5936 => x"76",     5937 => x"74",     5938 => x"71",     5939 => x"73",     5940 => x"76",     5941 => x"79",     5942 => x"77",     5943 => x"76", 
    5944 => x"74",     5945 => x"75",     5946 => x"7A",     5947 => x"79",     5948 => x"7A",     5949 => x"78",     5950 => x"79",     5951 => x"79", 
    5952 => x"7B",     5953 => x"7B",     5954 => x"77",     5955 => x"7A",     5956 => x"75",     5957 => x"78",     5958 => x"75",     5959 => x"77", 
    5960 => x"74",     5961 => x"78",     5962 => x"79",     5963 => x"74",     5964 => x"74",     5965 => x"72",     5966 => x"74",     5967 => x"76", 
    5968 => x"76",     5969 => x"73",     5970 => x"73",     5971 => x"74",     5972 => x"76",     5973 => x"7A",     5974 => x"77",     5975 => x"77", 
    5976 => x"77",     5977 => x"79",     5978 => x"7B",     5979 => x"78",     5980 => x"77",     5981 => x"75",     5982 => x"79",     5983 => x"78", 
    5984 => x"79",     5985 => x"77",     5986 => x"77",     5987 => x"79",     5988 => x"79",     5989 => x"79",     5990 => x"79",     5991 => x"7B", 
    5992 => x"77",     5993 => x"78",     5994 => x"72",     5995 => x"71",     5996 => x"70",     5997 => x"74",     5998 => x"75",     5999 => x"74", 
    6000 => x"72",     6001 => x"71",     6002 => x"75",     6003 => x"78",     6004 => x"7C",     6005 => x"77",     6006 => x"78",     6007 => x"78", 
    6008 => x"7A",     6009 => x"7A",     6010 => x"78",     6011 => x"78",     6012 => x"76",     6013 => x"7A",     6014 => x"76",     6015 => x"78", 
    6016 => x"75",     6017 => x"76",     6018 => x"77",     6019 => x"77",     6020 => x"78",     6021 => x"74",     6022 => x"76",     6023 => x"73", 
    6024 => x"76",     6025 => x"74",     6026 => x"77",     6027 => x"74",     6028 => x"75",     6029 => x"72",     6030 => x"74",     6031 => x"73", 
    6032 => x"73",     6033 => x"76",     6034 => x"71",     6035 => x"73",     6036 => x"74",     6037 => x"77",     6038 => x"78",     6039 => x"77", 
    6040 => x"76",     6041 => x"77",     6042 => x"7B",     6043 => x"7B",     6044 => x"7D",     6045 => x"77",     6046 => x"77",     6047 => x"75", 
    6048 => x"78",     6049 => x"76",     6050 => x"75",     6051 => x"75",     6052 => x"73",     6053 => x"76",     6054 => x"74",     6055 => x"75", 
    6056 => x"74",     6057 => x"76",     6058 => x"75",     6059 => x"74",     6060 => x"73",     6061 => x"73",     6062 => x"74",     6063 => x"73", 
    6064 => x"75",     6065 => x"73",     6066 => x"75",     6067 => x"75",     6068 => x"76",     6069 => x"75",     6070 => x"75",     6071 => x"77", 
    6072 => x"77",     6073 => x"7A",     6074 => x"78",     6075 => x"79",     6076 => x"76",     6077 => x"7B",     6078 => x"79",     6079 => x"77", 
    6080 => x"75",     6081 => x"72",     6082 => x"73",     6083 => x"73",     6084 => x"71",     6085 => x"71",     6086 => x"73",     6087 => x"73", 
    6088 => x"76",     6089 => x"75",     6090 => x"76",     6091 => x"75",     6092 => x"77",     6093 => x"77",     6094 => x"76",     6095 => x"77", 
    6096 => x"73",     6097 => x"76",     6098 => x"75",     6099 => x"76",     6100 => x"75",     6101 => x"74",     6102 => x"77",     6103 => x"78", 
    6104 => x"79",     6105 => x"78",     6106 => x"78",     6107 => x"77",     6108 => x"7C",     6109 => x"78",     6110 => x"77",     6111 => x"77", 
    6112 => x"75",     6113 => x"78",     6114 => x"76",     6115 => x"74",     6116 => x"72",     6117 => x"72",     6118 => x"74",     6119 => x"75", 
    6120 => x"74",     6121 => x"73",     6122 => x"74",     6123 => x"77",     6124 => x"79",     6125 => x"78",     6126 => x"75",     6127 => x"75", 
    6128 => x"79",     6129 => x"79",     6130 => x"77",     6131 => x"77",     6132 => x"74",     6133 => x"79",     6134 => x"78",     6135 => x"7A", 
    6136 => x"78",     6137 => x"77",     6138 => x"77",     6139 => x"77",     6140 => x"76",     6141 => x"77",     6142 => x"77",     6143 => x"78", 
    6144 => x"78",     6145 => x"76",     6146 => x"78",     6147 => x"73",     6148 => x"75",     6149 => x"76",     6150 => x"76",     6151 => x"75", 
    6152 => x"75",     6153 => x"74",     6154 => x"77",     6155 => x"77",     6156 => x"76",     6157 => x"75",     6158 => x"77",     6159 => x"79", 
    6160 => x"78",     6161 => x"79",     6162 => x"76",     6163 => x"78",     6164 => x"79",     6165 => x"78",     6166 => x"77",     6167 => x"76", 
    6168 => x"75",     6169 => x"77",     6170 => x"77",     6171 => x"75",     6172 => x"73",     6173 => x"74",     6174 => x"76",     6175 => x"77", 
    6176 => x"75",     6177 => x"75",     6178 => x"75",     6179 => x"79",     6180 => x"75",     6181 => x"75",     6182 => x"73",     6183 => x"74", 
    6184 => x"76",     6185 => x"77",     6186 => x"75",     6187 => x"74",     6188 => x"76",     6189 => x"76",     6190 => x"79",     6191 => x"78", 
    6192 => x"77",     6193 => x"76",     6194 => x"77",     6195 => x"77",     6196 => x"78",     6197 => x"76",     6198 => x"75",     6199 => x"76", 
    6200 => x"76",     6201 => x"77",     6202 => x"75",     6203 => x"74",     6204 => x"75",     6205 => x"76",     6206 => x"77",     6207 => x"78", 
    6208 => x"75",     6209 => x"76",     6210 => x"76",     6211 => x"76",     6212 => x"76",     6213 => x"75",     6214 => x"76",     6215 => x"76", 
    6216 => x"77",     6217 => x"78",     6218 => x"76",     6219 => x"77",     6220 => x"77",     6221 => x"77",     6222 => x"76",     6223 => x"74", 
    6224 => x"75",     6225 => x"76",     6226 => x"76",     6227 => x"74",     6228 => x"75",     6229 => x"74",     6230 => x"77",     6231 => x"76", 
    6232 => x"75",     6233 => x"76",     6234 => x"77",     6235 => x"78",     6236 => x"79",     6237 => x"77",     6238 => x"74",     6239 => x"76", 
    6240 => x"74",     6241 => x"75",     6242 => x"75",     6243 => x"75",     6244 => x"75",     6245 => x"75",     6246 => x"76",     6247 => x"77", 
    6248 => x"78",     6249 => x"77",     6250 => x"79",     6251 => x"77",     6252 => x"76",     6253 => x"76",     6254 => x"76",     6255 => x"77", 
    6256 => x"74",     6257 => x"75",     6258 => x"73",     6259 => x"76",     6260 => x"75",     6261 => x"77",     6262 => x"75",     6263 => x"77", 
    6264 => x"77",     6265 => x"77",     6266 => x"77",     6267 => x"75",     6268 => x"75",     6269 => x"74",     6270 => x"74",     6271 => x"75", 
    6272 => x"76",     6273 => x"75",     6274 => x"77",     6275 => x"77",     6276 => x"78",     6277 => x"77",     6278 => x"76",     6279 => x"76", 
    6280 => x"77",     6281 => x"76",     6282 => x"75",     6283 => x"76",     6284 => x"76",     6285 => x"77",     6286 => x"78",     6287 => x"76", 
    6288 => x"76",     6289 => x"76",     6290 => x"76",     6291 => x"76",     6292 => x"76",     6293 => x"76",     6294 => x"75",     6295 => x"78", 
    6296 => x"76",     6297 => x"77",     6298 => x"78",     6299 => x"78",     6300 => x"77",     6301 => x"76",     6302 => x"76",     6303 => x"77", 
    6304 => x"78",     6305 => x"76",     6306 => x"75",     6307 => x"75",     6308 => x"76",     6309 => x"77",     6310 => x"77",     6311 => x"74", 
    6312 => x"76",     6313 => x"76",     6314 => x"78",     6315 => x"77",     6316 => x"76",     6317 => x"75",     6318 => x"76",     6319 => x"76", 
    6320 => x"77",     6321 => x"74",     6322 => x"76",     6323 => x"75",     6324 => x"76",     6325 => x"77",     6326 => x"77",     6327 => x"77", 
    6328 => x"76",     6329 => x"76",     6330 => x"76",     6331 => x"76",     6332 => x"75",     6333 => x"75",     6334 => x"75",     6335 => x"78", 
    6336 => x"76",     6337 => x"78",     6338 => x"76",     6339 => x"76",     6340 => x"77",     6341 => x"78",     6342 => x"77",     6343 => x"76", 
    6344 => x"76",     6345 => x"75",     6346 => x"76",     6347 => x"74",     6348 => x"76",     6349 => x"76",     6350 => x"75",     6351 => x"74", 
    6352 => x"74",     6353 => x"76",     6354 => x"76",     6355 => x"78",     6356 => x"76",     6357 => x"75",     6358 => x"75",     6359 => x"76", 
    6360 => x"76",     6361 => x"76",     6362 => x"76",     6363 => x"75",     6364 => x"78",     6365 => x"77",     6366 => x"76",     6367 => x"76", 
    6368 => x"76",     6369 => x"78",     6370 => x"77",     6371 => x"78",     6372 => x"75",     6373 => x"77",     6374 => x"76",     6375 => x"76", 
    6376 => x"76",     6377 => x"75",     6378 => x"77",     6379 => x"77",     6380 => x"76",     6381 => x"74",     6382 => x"75",     6383 => x"74", 
    6384 => x"77",     6385 => x"76",     6386 => x"77",     6387 => x"75",     6388 => x"76",     6389 => x"76",     6390 => x"77",     6391 => x"76", 
    6392 => x"75",     6393 => x"76",     6394 => x"75",     6395 => x"78",     6396 => x"76",     6397 => x"76",     6398 => x"75",     6399 => x"76", 
    6400 => x"77",     6401 => x"77",     6402 => x"77",     6403 => x"77",     6404 => x"78",     6405 => x"77",     6406 => x"78",     6407 => x"77", 
    6408 => x"77",     6409 => x"77",     6410 => x"77",     6411 => x"76",     6412 => x"75",     6413 => x"75",     6414 => x"76",     6415 => x"76", 
    6416 => x"75",     6417 => x"75",     6418 => x"74",     6419 => x"76",     6420 => x"75",     6421 => x"77",     6422 => x"77",     6423 => x"76", 
    6424 => x"78",     6425 => x"77",     6426 => x"78",     6427 => x"76",     6428 => x"76",     6429 => x"75",     6430 => x"77"
);


    --constant sLUT : sine_table_t := (
    --    0 => x"80",  1 => x"86",  2 => x"8C",  3 => x"92",
    --    4 => x"98",  5 => x"9E",  6 => x"A5",  7 => x"AA",
    --    8 => x"B0",  9 => x"B6", 10 => x"BC", 11 => x"C1",
    --    12 => x"C6", 13 => x"CB", 14 => x"D0", 15 => x"D5",
    --    16 => x"DA", 17 => x"DE", 18 => x"E2", 19 => x"E6",
    --    20 => x"EA", 21 => x"ED", 22 => x"F0", 23 => x"F3",
    --    24 => x"F5", 25 => x"F8", 26 => x"FA", 27 => x"FB",
    --    28 => x"FD", 29 => x"FE", 30 => x"FE", 31 => x"FF",
    --    32 => x"FF", 33 => x"FF", 34 => x"FE", 35 => x"FE",
    --    36 => x"FD", 37 => x"FB", 38 => x"FA", 39 => x"F8",
    --    40 => x"F5", 41 => x"F3", 42 => x"F0", 43 => x"ED",
    --    44 => x"EA", 45 => x"E6", 46 => x"E2", 47 => x"DE",
    --    48 => x"DA", 49 => x"D5", 50 => x"D0", 51 => x"CB",
    --    52 => x"C6", 53 => x"C1", 54 => x"BC", 55 => x"B6",
    --    56 => x"B0", 57 => x"AA", 58 => x"A5", 59 => x"9E",
    --    60 => x"98", 61 => x"92", 62 => x"8C", 63 => x"86",
    --    64 => x"80", 65 => x"79", 66 => x"73", 67 => x"6D",
    --    68 => x"67", 69 => x"61", 70 => x"5A", 71 => x"55",
    --    72 => x"4F", 73 => x"49", 74 => x"43", 75 => x"3E",
    --    76 => x"39", 77 => x"34", 78 => x"2F", 79 => x"2A",
    --    80 => x"25", 81 => x"21", 82 => x"1D", 83 => x"19",
    --    84 => x"15", 85 => x"12", 86 => x"0F", 87 => x"0C",
    --    88 => x"0A", 89 => x"07", 90 => x"05", 91 => x"04",
    --    92 => x"02", 93 => x"01", 94 => x"01", 95 => x"00",
    --    96 => x"00", 97 => x"00", 98 => x"01", 99 => x"01",
    --    100 => x"02",101 => x"04",102 => x"05",103 => x"07",
    --    104 => x"0A",105 => x"0C",106 => x"0F",107 => x"12",
    --    108 => x"15",109 => x"19",110 => x"1D",111 => x"21",
    --    112 => x"25",113 => x"2A",114 => x"2F",115 => x"34",
    --    116 => x"39",117 => x"3E",118 => x"43",119 => x"49",
    --    120 => x"4F",121 => x"55",122 => x"5A",123 => x"61",
    --    124 => x"67",125 => x"6D",126 => x"73",127 => x"79"
    --);



    signal vwoop_sig : std_logic_vector(7 downto 0); 
    signal snake_sig : std_logic_vector(7 downto 0);
    signal womps_sig : std_logic_vector(7 downto 0); 

    signal vwoop_going  : std_logic; 
    signal liz_going    : std_logic; 
    signal womp_going   : std_logic;

    signal audio_cnt_1   : integer; 
    signal audio_cnt_2   : integer; 
    signal audio_cnt_3   : integer; 

    signal clk_div_cnt_1 : integer;
    signal clk_div_cnt_2 : integer;
    signal clk_div_cnt_3 : integer;

    signal audio_cnt   : integer; 

    signal clk_div_cnt : integer;

    signal twisty_turn_d  : std_logic := '0';
signal chompy_appy_d  : std_logic := '0';

begin 

    --chompy_appy : in  std_logic; 
    --twisty_turn : in  std_logic; 
    --ha_loser    : in  std_logic; 
   
vwoop_sound : process(clk, rst)
begin
    if rst = '1' then
        audio_cnt_1    <= 0;
        clk_div_cnt_1  <= 0;
        vwoop_going    <= '0';
        vwoop_sig      <= (others => '0');
        twisty_turn_d  <= '0';

    elsif rising_edge(clk) then

        -- Edge detect
        twisty_turn_d <= twisty_turn;

        if twisty_turn = '1' and twisty_turn_d = '0' then
            vwoop_going   <= '1';
            audio_cnt_1   <= 0;
            clk_div_cnt_1 <= 0;
        end if;

        -- Divider
        if clk_div_cnt_1 = 6249 then
            clk_div_cnt_1 <= 0;

            if vwoop_going = '1' then
                vwoop_sig <= vwoopLUT(audio_cnt_1);

                if audio_cnt_1 = vwoop_len-1 then
                    audio_cnt_1 <= 0;
                    vwoop_going <= '0';
                else
                    audio_cnt_1 <= audio_cnt_1 + 1;
                end if;
            end if;

        else
            clk_div_cnt_1 <= clk_div_cnt_1 + 1;
        end if;

    end if;
end process;

snake_sound : process(clk, rst)
begin
    if rst = '1' then
        audio_cnt_2    <= 0;
        clk_div_cnt_2  <= 0;
        liz_going      <= '0';
        snake_sig      <= (others => '0');
        chompy_appy_d  <= '0';

    elsif rising_edge(clk) then

        -- Edge detect
        chompy_appy_d <= chompy_appy;

        if chompy_appy = '1' and chompy_appy_d = '0' then
            liz_going     <= '1';
            audio_cnt_2   <= 0;
            clk_div_cnt_2 <= 0;
        end if;

        if clk_div_cnt_2 = 6249 then
            clk_div_cnt_2 <= 0;

            if liz_going = '1' then
                snake_sig <= lizLUT(audio_cnt_2);

                if audio_cnt_2 = liz_len-1 then
                    audio_cnt_2 <= 0;
                    liz_going   <= '0';
                else
                    audio_cnt_2 <= audio_cnt_2 + 1;
                end if;
            end if;

        else
            clk_div_cnt_2 <= clk_div_cnt_2 + 1;
        end if;

    end if;
end process;

womp_sound : process(clk, rst)
begin
    if rst = '1' then
        audio_cnt_3    <= 0;
        clk_div_cnt_3  <= 0;
        womp_going     <= '0';
        womps_sig      <= (others => '0');

    elsif rising_edge(clk) then

        -- reuse chompy_appy_d from snake process
        if chompy_appy = '1' and chompy_appy_d = '0' then
            womp_going    <= '1';
            audio_cnt_3   <= 0;
            clk_div_cnt_3 <= 0;
        end if;

        if clk_div_cnt_3 = 6249 then
            clk_div_cnt_3 <= 0;

            if womp_going = '1' then
                womps_sig <= wompLUT(audio_cnt_3);

                if audio_cnt_3 = womp_len-1 then
                    audio_cnt_3 <= 0;
                    womp_going  <= '0';
                else
                    audio_cnt_3 <= audio_cnt_3 + 1;
                end if;
            end if;

        else
            clk_div_cnt_3 <= clk_div_cnt_3 + 1;
        end if;

    end if;
end process;

audio_mux : process(clk, rst)
begin
    if rst = '1' then
        audio_out <= (others => '0');

    elsif rising_edge(clk) then

        audio_out <= (others => '0');

        if vwoop_going = '1' then
            audio_out <= vwoop_sig;
        end if;

        if liz_going = '1' then
            audio_out <= snake_sig;
        end if;

        if womp_going = '1' then
            audio_out <= womps_sig;
        end if;

    end if;
end process;
   
--    vwoop_sound : process(clk, rst) is begin
--        if rst = '1' then
--            audio_cnt_1 <= 0;
--            clk_div_cnt_1 <= 0; 
--            vwoop_going <= '0';
--        elsif rising_edge(clk) then
--            if twisty_turn = '1' then 
--                vwoop_going <= '1';
--                audio_cnt_1 <= 0;
--                clk_div_cnt_1 <= 0; 
--            end if; 
--            clk_div_cnt_1 <= clk_div_cnt_1 + 1;
--            if clk_div_cnt_1 = 6250 then 
--                clk_div_cnt_1 <= 0;
--                vwoop_sig <= vwoopLUT(audio_cnt_1); 
--   
--                audio_cnt_1 <= audio_cnt_1 + 1; 
--   
--                if audio_cnt_1 = vwoop_len then
--                    audio_cnt_1 <= 0; 
--                    vwoop_going <= '0';
--                end if; 
--            end if; 
--        end if; 
--    end process vwoop_sound; 
--   
--    snake_sound : process(clk, rst) is begin
--        if rst = '1' then
--            audio_cnt_2 <= 0;
--            clk_div_cnt_2 <= 0; 
--            liz_going <= '0';
--        elsif rising_edge(clk) then
--            if chompy_appy = '1' then 
--                liz_going <= '1';
--                audio_cnt_2 <= 0;
--                clk_div_cnt_2 <= 0; 
--            end if; 
--            clk_div_cnt_2 <= clk_div_cnt_2 + 1;
--            if clk_div_cnt_2 = 6250 then 
--                clk_div_cnt_2 <= 0;
--                snake_sig <= lizLUT(audio_cnt_2); 
--   
--                audio_cnt_2 <= audio_cnt_2 + 1; 
--   
--                if audio_cnt_2 = liz_len then
--                    audio_cnt_2 <= 0; 
--                    liz_going <= '0';
--                end if; 
--            end if; 
--        end if; 
--    end process snake_sound; 
--   
--    womp_sound : process(clk, rst) is begin
--        if rst = '1' then
--            audio_cnt_3 <= 0;
--            clk_div_cnt_3 <= 0; 
--            womp_going <= '0';
--        elsif rising_edge(clk) then
--            if chompy_appy = '1' then 
--                womp_going <= '1';
--                audio_cnt_3 <= 0;
--                clk_div_cnt_3 <= 0; 
--            end if; 
--            clk_div_cnt_3 <= clk_div_cnt_3 + 1;
--            if clk_div_cnt_3 = 6250 then 
--                clk_div_cnt_3 <= 0;
--                womps_sig <= wompLUT(audio_cnt_3); 
--   
--                audio_cnt_3 <= audio_cnt_3 + 1; 
--   
--                if audio_cnt_3 = womp_len then
--                    audio_cnt_3 <= 0; 
--                    womp_going <= '0';
--                end if; 
--            end if; 
--        end if; 
--    end process womp_sound; 
--   
--   audio_mux : process(clk, rst) is begin 
--    if rst = '1' then
--        audio_out <= (others => '0'); 
--    elsif rising_edge(clk) then
--        audio_out <= (others => '0'); 
--        if vwoop_going = '1' then
--            audio_out <= vwoop_sig; 
--        end if; 
--        if liz_going = '1' then 
--            audio_out <= snake_sig; 
--        end if; 
--        if womp_going = '1' then 
--            audio_out <= womps_sig; 
--        end if;
--    end if; 
--   end process audio_mux; 

--    sfx : process(clk, rst) is begin 
--        if rst = '1' then 
--            audio_out   <= (others => '0');
--
--            clk_div_cnt <= 0; 
--            audio_cnt   <= 0; 
--        elsif rising_edge(clk) then 
--            if clk_div_cnt = 6250 then
--                if audio_cnt < liz_len then 
--                    audio_out <= lizLUT(audio_cnt);
--
--                elsif audio_cnt < liz_len + womp_len then
--                    audio_out <= wompLUT(audio_cnt - liz_len);
--
--                else
--                    audio_out <= vwoopLUT(audio_cnt - liz_len - womp_len);
--                end if;
--                            
--                audio_cnt <= audio_cnt + 1; 
--
--                if audio_cnt >= liz_len + womp_len + vwoop_len then
--                    audio_cnt <= 0; 
--                end if; 
--
--                clk_div_cnt <= 0; 
--            else
--                clk_div_cnt <= clk_div_cnt + 1; 
--            end if;      
--        end if; 
--    end process sfx; 
--
end architecture arch; 

